// amm_master_qsys_custom_with_bfm_tb.v

// Generated using ACDS version 13.0sp1 232 at 2015.02.16.16:52:33

`timescale 1 ps / 1 ps
module amm_master_qsys_custom_with_bfm_tb (
	);

	wire    amm_master_qsys_custom_with_bfm_inst_clk_bfm_clk_clk;       // amm_master_qsys_custom_with_bfm_inst_clk_bfm:clk -> [amm_master_qsys_custom_with_bfm_inst:clk_clk, amm_master_qsys_custom_with_bfm_inst_reset_bfm:clk]
	wire    amm_master_qsys_custom_with_bfm_inst_reset_bfm_reset_reset; // amm_master_qsys_custom_with_bfm_inst_reset_bfm:reset -> amm_master_qsys_custom_with_bfm_inst:reset_reset_n

	amm_master_qsys_custom_with_bfm amm_master_qsys_custom_with_bfm_inst (
		.clk_clk                            (amm_master_qsys_custom_with_bfm_inst_clk_bfm_clk_clk),       //                   clk.clk
		.reset_reset_n                      (amm_master_qsys_custom_with_bfm_inst_reset_bfm_reset_reset), //                 reset.reset_n
		.custom_module_conduit_rdwr_cntl    (),                                                           // custom_module_conduit.rdwr_cntl
		.custom_module_conduit_n_action     (),                                                           //                      .n_action
		.custom_module_conduit_add_data_sel (),                                                           //                      .add_data_sel
		.custom_module_conduit_rdwr_address ()                                                            //                      .rdwr_address
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) amm_master_qsys_custom_with_bfm_inst_clk_bfm (
		.clk (amm_master_qsys_custom_with_bfm_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) amm_master_qsys_custom_with_bfm_inst_reset_bfm (
		.reset (amm_master_qsys_custom_with_bfm_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (amm_master_qsys_custom_with_bfm_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
