// amm_master_qsys.v

// Generated using ACDS version 13.0sp1 232 at 2014.11.03.12:20:42

`timescale 1 ps / 1 ps
module amm_master_qsys (
		input  wire        clk_clk,                             //                         clk.clk
		input  wire        reset_reset_n,                       //                       reset.reset_n
		output wire [11:0] new_sdram_controller_0_wire_addr,    // new_sdram_controller_0_wire.addr
		output wire [1:0]  new_sdram_controller_0_wire_ba,      //                            .ba
		output wire        new_sdram_controller_0_wire_cas_n,   //                            .cas_n
		output wire        new_sdram_controller_0_wire_cke,     //                            .cke
		output wire        new_sdram_controller_0_wire_cs_n,    //                            .cs_n
		inout  wire [31:0] new_sdram_controller_0_wire_dq,      //                            .dq
		output wire [3:0]  new_sdram_controller_0_wire_dqm,     //                            .dqm
		output wire        new_sdram_controller_0_wire_ras_n,   //                            .ras_n
		output wire        new_sdram_controller_0_wire_we_n,    //                            .we_n
		input  wire        write_master_control_fixed_location, //        write_master_control.fixed_location
		input  wire [25:0] write_master_control_write_base,     //                            .write_base
		input  wire [25:0] write_master_control_write_length,   //                            .write_length
		input  wire        write_master_control_go,             //                            .go
		output wire        write_master_control_done,           //                            .done
		input  wire        write_master_user_write_buffer,      //           write_master_user.write_buffer
		input  wire [31:0] write_master_user_buffer_input_data, //                            .buffer_input_data
		output wire        write_master_user_buffer_full,       //                            .buffer_full
		input  wire        read_master_control_fixed_location,  //         read_master_control.fixed_location
		input  wire [25:0] read_master_control_read_base,       //                            .read_base
		input  wire [25:0] read_master_control_read_length,     //                            .read_length
		input  wire        read_master_control_go,              //                            .go
		output wire        read_master_control_done,            //                            .done
		output wire        read_master_control_early_done,      //                            .early_done
		input  wire        read_master_user_read_buffer,        //            read_master_user.read_buffer
		output wire [31:0] read_master_user_buffer_output_data, //                            .buffer_output_data
		output wire        read_master_user_data_available      //                            .data_available
	);

	wire         write_master_avalon_master_waitrequest;                                                         // write_master_avalon_master_translator:av_waitrequest -> write_master:master_waitrequest
	wire  [31:0] write_master_avalon_master_writedata;                                                           // write_master:master_writedata -> write_master_avalon_master_translator:av_writedata
	wire  [25:0] write_master_avalon_master_address;                                                             // write_master:master_address -> write_master_avalon_master_translator:av_address
	wire         write_master_avalon_master_write;                                                               // write_master:master_write -> write_master_avalon_master_translator:av_write
	wire   [3:0] write_master_avalon_master_byteenable;                                                          // write_master:master_byteenable -> write_master_avalon_master_translator:av_byteenable
	wire         read_master_avalon_master_waitrequest;                                                          // read_master_avalon_master_translator:av_waitrequest -> read_master:master_waitrequest
	wire  [25:0] read_master_avalon_master_address;                                                              // read_master:master_address -> read_master_avalon_master_translator:av_address
	wire         read_master_avalon_master_read;                                                                 // read_master:master_read -> read_master_avalon_master_translator:av_read
	wire  [31:0] read_master_avalon_master_readdata;                                                             // read_master_avalon_master_translator:av_readdata -> read_master:master_readdata
	wire         read_master_avalon_master_readdatavalid;                                                        // read_master_avalon_master_translator:av_readdatavalid -> read_master:master_readdatavalid
	wire   [3:0] read_master_avalon_master_byteenable;                                                           // read_master:master_byteenable -> read_master_avalon_master_translator:av_byteenable
	wire         new_sdram_controller_0_s1_translator_avalon_anti_slave_0_waitrequest;                           // new_sdram_controller_0:za_waitrequest -> new_sdram_controller_0_s1_translator:av_waitrequest
	wire  [31:0] new_sdram_controller_0_s1_translator_avalon_anti_slave_0_writedata;                             // new_sdram_controller_0_s1_translator:av_writedata -> new_sdram_controller_0:az_data
	wire  [23:0] new_sdram_controller_0_s1_translator_avalon_anti_slave_0_address;                               // new_sdram_controller_0_s1_translator:av_address -> new_sdram_controller_0:az_addr
	wire         new_sdram_controller_0_s1_translator_avalon_anti_slave_0_chipselect;                            // new_sdram_controller_0_s1_translator:av_chipselect -> new_sdram_controller_0:az_cs
	wire         new_sdram_controller_0_s1_translator_avalon_anti_slave_0_write;                                 // new_sdram_controller_0_s1_translator:av_write -> new_sdram_controller_0:az_wr_n
	wire         new_sdram_controller_0_s1_translator_avalon_anti_slave_0_read;                                  // new_sdram_controller_0_s1_translator:av_read -> new_sdram_controller_0:az_rd_n
	wire  [31:0] new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdata;                              // new_sdram_controller_0:za_data -> new_sdram_controller_0_s1_translator:av_readdata
	wire         new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdatavalid;                         // new_sdram_controller_0:za_valid -> new_sdram_controller_0_s1_translator:av_readdatavalid
	wire   [3:0] new_sdram_controller_0_s1_translator_avalon_anti_slave_0_byteenable;                            // new_sdram_controller_0_s1_translator:av_byteenable -> new_sdram_controller_0:az_be_n
	wire         write_master_avalon_master_translator_avalon_universal_master_0_waitrequest;                    // write_master_avalon_master_translator_avalon_universal_master_0_agent:av_waitrequest -> write_master_avalon_master_translator:uav_waitrequest
	wire   [2:0] write_master_avalon_master_translator_avalon_universal_master_0_burstcount;                     // write_master_avalon_master_translator:uav_burstcount -> write_master_avalon_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] write_master_avalon_master_translator_avalon_universal_master_0_writedata;                      // write_master_avalon_master_translator:uav_writedata -> write_master_avalon_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [25:0] write_master_avalon_master_translator_avalon_universal_master_0_address;                        // write_master_avalon_master_translator:uav_address -> write_master_avalon_master_translator_avalon_universal_master_0_agent:av_address
	wire         write_master_avalon_master_translator_avalon_universal_master_0_lock;                           // write_master_avalon_master_translator:uav_lock -> write_master_avalon_master_translator_avalon_universal_master_0_agent:av_lock
	wire         write_master_avalon_master_translator_avalon_universal_master_0_write;                          // write_master_avalon_master_translator:uav_write -> write_master_avalon_master_translator_avalon_universal_master_0_agent:av_write
	wire         write_master_avalon_master_translator_avalon_universal_master_0_read;                           // write_master_avalon_master_translator:uav_read -> write_master_avalon_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] write_master_avalon_master_translator_avalon_universal_master_0_readdata;                       // write_master_avalon_master_translator_avalon_universal_master_0_agent:av_readdata -> write_master_avalon_master_translator:uav_readdata
	wire         write_master_avalon_master_translator_avalon_universal_master_0_debugaccess;                    // write_master_avalon_master_translator:uav_debugaccess -> write_master_avalon_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] write_master_avalon_master_translator_avalon_universal_master_0_byteenable;                     // write_master_avalon_master_translator:uav_byteenable -> write_master_avalon_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         write_master_avalon_master_translator_avalon_universal_master_0_readdatavalid;                  // write_master_avalon_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> write_master_avalon_master_translator:uav_readdatavalid
	wire         read_master_avalon_master_translator_avalon_universal_master_0_waitrequest;                     // read_master_avalon_master_translator_avalon_universal_master_0_agent:av_waitrequest -> read_master_avalon_master_translator:uav_waitrequest
	wire   [2:0] read_master_avalon_master_translator_avalon_universal_master_0_burstcount;                      // read_master_avalon_master_translator:uav_burstcount -> read_master_avalon_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] read_master_avalon_master_translator_avalon_universal_master_0_writedata;                       // read_master_avalon_master_translator:uav_writedata -> read_master_avalon_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [25:0] read_master_avalon_master_translator_avalon_universal_master_0_address;                         // read_master_avalon_master_translator:uav_address -> read_master_avalon_master_translator_avalon_universal_master_0_agent:av_address
	wire         read_master_avalon_master_translator_avalon_universal_master_0_lock;                            // read_master_avalon_master_translator:uav_lock -> read_master_avalon_master_translator_avalon_universal_master_0_agent:av_lock
	wire         read_master_avalon_master_translator_avalon_universal_master_0_write;                           // read_master_avalon_master_translator:uav_write -> read_master_avalon_master_translator_avalon_universal_master_0_agent:av_write
	wire         read_master_avalon_master_translator_avalon_universal_master_0_read;                            // read_master_avalon_master_translator:uav_read -> read_master_avalon_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] read_master_avalon_master_translator_avalon_universal_master_0_readdata;                        // read_master_avalon_master_translator_avalon_universal_master_0_agent:av_readdata -> read_master_avalon_master_translator:uav_readdata
	wire         read_master_avalon_master_translator_avalon_universal_master_0_debugaccess;                     // read_master_avalon_master_translator:uav_debugaccess -> read_master_avalon_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] read_master_avalon_master_translator_avalon_universal_master_0_byteenable;                      // read_master_avalon_master_translator:uav_byteenable -> read_master_avalon_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         read_master_avalon_master_translator_avalon_universal_master_0_readdatavalid;                   // read_master_avalon_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> read_master_avalon_master_translator:uav_readdatavalid
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // new_sdram_controller_0_s1_translator:uav_waitrequest -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;              // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> new_sdram_controller_0_s1_translator:uav_burstcount
	wire  [31:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;               // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> new_sdram_controller_0_s1_translator:uav_writedata
	wire  [25:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                 // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> new_sdram_controller_0_s1_translator:uav_address
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                   // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> new_sdram_controller_0_s1_translator:uav_write
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                    // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> new_sdram_controller_0_s1_translator:uav_lock
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                    // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> new_sdram_controller_0_s1_translator:uav_read
	wire  [31:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                // new_sdram_controller_0_s1_translator:uav_readdata -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // new_sdram_controller_0_s1_translator:uav_readdatavalid -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> new_sdram_controller_0_s1_translator:uav_debugaccess
	wire   [3:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;              // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> new_sdram_controller_0_s1_translator:uav_byteenable
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;            // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [93:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;             // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;            // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [93:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         write_master_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket;           // write_master_avalon_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         write_master_avalon_master_translator_avalon_universal_master_0_agent_cp_valid;                 // write_master_avalon_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         write_master_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket;         // write_master_avalon_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [92:0] write_master_avalon_master_translator_avalon_universal_master_0_agent_cp_data;                  // write_master_avalon_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         write_master_avalon_master_translator_avalon_universal_master_0_agent_cp_ready;                 // addr_router:sink_ready -> write_master_avalon_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         read_master_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket;            // read_master_avalon_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         read_master_avalon_master_translator_avalon_universal_master_0_agent_cp_valid;                  // read_master_avalon_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         read_master_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket;          // read_master_avalon_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [92:0] read_master_avalon_master_translator_avalon_universal_master_0_agent_cp_data;                   // read_master_avalon_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         read_master_avalon_master_translator_avalon_universal_master_0_agent_cp_ready;                  // addr_router_001:sink_ready -> read_master_avalon_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                   // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [92:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                    // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router:sink_ready -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         rst_controller_reset_out_reset;                                                                 // rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, id_router:reset, new_sdram_controller_0:reset_n, new_sdram_controller_0_s1_translator:reset, new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:reset, new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, read_master:reset, read_master_avalon_master_translator:reset, read_master_avalon_master_translator_avalon_universal_master_0_agent:reset, rsp_xbar_demux:reset, write_master:reset, write_master_avalon_master_translator:reset, write_master_avalon_master_translator_avalon_universal_master_0_agent:reset]
	wire         cmd_xbar_demux_src0_endofpacket;                                                                // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                      // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                              // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [92:0] cmd_xbar_demux_src0_data;                                                                       // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [1:0] cmd_xbar_demux_src0_channel;                                                                    // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                      // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                            // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                  // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                          // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [92:0] cmd_xbar_demux_001_src0_data;                                                                   // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [1:0] cmd_xbar_demux_001_src0_channel;                                                                // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                  // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_src0_endofpacket;                                                                // rsp_xbar_demux:src0_endofpacket -> write_master_avalon_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                      // rsp_xbar_demux:src0_valid -> write_master_avalon_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                              // rsp_xbar_demux:src0_startofpacket -> write_master_avalon_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [92:0] rsp_xbar_demux_src0_data;                                                                       // rsp_xbar_demux:src0_data -> write_master_avalon_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [1:0] rsp_xbar_demux_src0_channel;                                                                    // rsp_xbar_demux:src0_channel -> write_master_avalon_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_demux_src1_endofpacket;                                                                // rsp_xbar_demux:src1_endofpacket -> read_master_avalon_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                      // rsp_xbar_demux:src1_valid -> read_master_avalon_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                              // rsp_xbar_demux:src1_startofpacket -> read_master_avalon_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [92:0] rsp_xbar_demux_src1_data;                                                                       // rsp_xbar_demux:src1_data -> read_master_avalon_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [1:0] rsp_xbar_demux_src1_channel;                                                                    // rsp_xbar_demux:src1_channel -> read_master_avalon_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         addr_router_src_endofpacket;                                                                    // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         addr_router_src_valid;                                                                          // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire         addr_router_src_startofpacket;                                                                  // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [92:0] addr_router_src_data;                                                                           // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire   [1:0] addr_router_src_channel;                                                                        // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire         addr_router_src_ready;                                                                          // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire         rsp_xbar_demux_src0_ready;                                                                      // write_master_avalon_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux:src0_ready
	wire         addr_router_001_src_endofpacket;                                                                // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         addr_router_001_src_valid;                                                                      // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire         addr_router_001_src_startofpacket;                                                              // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [92:0] addr_router_001_src_data;                                                                       // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire   [1:0] addr_router_001_src_channel;                                                                    // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire         addr_router_001_src_ready;                                                                      // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire         rsp_xbar_demux_src1_ready;                                                                      // read_master_avalon_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux:src1_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                   // cmd_xbar_mux:src_endofpacket -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                         // cmd_xbar_mux:src_valid -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                 // cmd_xbar_mux:src_startofpacket -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [92:0] cmd_xbar_mux_src_data;                                                                          // cmd_xbar_mux:src_data -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [1:0] cmd_xbar_mux_src_channel;                                                                       // cmd_xbar_mux:src_channel -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                         // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                      // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                            // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                    // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [92:0] id_router_src_data;                                                                             // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [1:0] id_router_src_channel;                                                                          // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                            // rsp_xbar_demux:sink_ready -> id_router:src_ready

	amm_master_qsys_new_sdram_controller_0 new_sdram_controller_0 (
		.clk            (clk_clk),                                                                //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                                        // reset.reset_n
		.az_addr        (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~new_sdram_controller_0_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~new_sdram_controller_0_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~new_sdram_controller_0_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (new_sdram_controller_0_wire_addr),                                       //  wire.export
		.zs_ba          (new_sdram_controller_0_wire_ba),                                         //      .export
		.zs_cas_n       (new_sdram_controller_0_wire_cas_n),                                      //      .export
		.zs_cke         (new_sdram_controller_0_wire_cke),                                        //      .export
		.zs_cs_n        (new_sdram_controller_0_wire_cs_n),                                       //      .export
		.zs_dq          (new_sdram_controller_0_wire_dq),                                         //      .export
		.zs_dqm         (new_sdram_controller_0_wire_dqm),                                        //      .export
		.zs_ras_n       (new_sdram_controller_0_wire_ras_n),                                      //      .export
		.zs_we_n        (new_sdram_controller_0_wire_we_n)                                        //      .export
	);

	custom_master #(
		.MASTER_DIRECTION    (1),
		.DATA_WIDTH          (32),
		.ADDRESS_WIDTH       (26),
		.BURST_CAPABLE       (0),
		.MAXIMUM_BURST_COUNT (2),
		.BURST_COUNT_WIDTH   (2),
		.FIFO_DEPTH          (16),
		.FIFO_DEPTH_LOG2     (4),
		.MEMORY_BASED_FIFO   (1)
	) write_master (
		.clk                     (clk_clk),                                //       clock_reset.clk
		.reset                   (rst_controller_reset_out_reset),         // clock_reset_reset.reset
		.master_address          (write_master_avalon_master_address),     //     avalon_master.address
		.master_write            (write_master_avalon_master_write),       //                  .write
		.master_byteenable       (write_master_avalon_master_byteenable),  //                  .byteenable
		.master_writedata        (write_master_avalon_master_writedata),   //                  .writedata
		.master_waitrequest      (write_master_avalon_master_waitrequest), //                  .waitrequest
		.control_fixed_location  (write_master_control_fixed_location),    //           control.export
		.control_write_base      (write_master_control_write_base),        //                  .export
		.control_write_length    (write_master_control_write_length),      //                  .export
		.control_go              (write_master_control_go),                //                  .export
		.control_done            (write_master_control_done),              //                  .export
		.user_write_buffer       (write_master_user_write_buffer),         //              user.export
		.user_buffer_input_data  (write_master_user_buffer_input_data),    //                  .export
		.user_buffer_full        (write_master_user_buffer_full),          //                  .export
		.master_read             (),                                       //       (terminated)
		.master_readdata         (32'b00000000000000000000000000000000),   //       (terminated)
		.master_readdatavalid    (1'b0),                                   //       (terminated)
		.master_burstcount       (),                                       //       (terminated)
		.control_read_base       (26'b00000000000000000000000000),         //       (terminated)
		.control_read_length     (26'b00000000000000000000000000),         //       (terminated)
		.control_early_done      (),                                       //       (terminated)
		.user_read_buffer        (1'b0),                                   //       (terminated)
		.user_buffer_output_data (),                                       //       (terminated)
		.user_data_available     ()                                        //       (terminated)
	);

	custom_master #(
		.MASTER_DIRECTION    (0),
		.DATA_WIDTH          (32),
		.ADDRESS_WIDTH       (26),
		.BURST_CAPABLE       (0),
		.MAXIMUM_BURST_COUNT (2),
		.BURST_COUNT_WIDTH   (2),
		.FIFO_DEPTH          (32),
		.FIFO_DEPTH_LOG2     (5),
		.MEMORY_BASED_FIFO   (1)
	) read_master (
		.clk                     (clk_clk),                                 //       clock_reset.clk
		.reset                   (rst_controller_reset_out_reset),          // clock_reset_reset.reset
		.master_address          (read_master_avalon_master_address),       //     avalon_master.address
		.master_read             (read_master_avalon_master_read),          //                  .read
		.master_byteenable       (read_master_avalon_master_byteenable),    //                  .byteenable
		.master_readdata         (read_master_avalon_master_readdata),      //                  .readdata
		.master_readdatavalid    (read_master_avalon_master_readdatavalid), //                  .readdatavalid
		.master_waitrequest      (read_master_avalon_master_waitrequest),   //                  .waitrequest
		.control_fixed_location  (read_master_control_fixed_location),      //           control.export
		.control_read_base       (read_master_control_read_base),           //                  .export
		.control_read_length     (read_master_control_read_length),         //                  .export
		.control_go              (read_master_control_go),                  //                  .export
		.control_done            (read_master_control_done),                //                  .export
		.control_early_done      (read_master_control_early_done),          //                  .export
		.user_read_buffer        (read_master_user_read_buffer),            //              user.export
		.user_buffer_output_data (read_master_user_buffer_output_data),     //                  .export
		.user_data_available     (read_master_user_data_available),         //                  .export
		.master_write            (),                                        //       (terminated)
		.master_writedata        (),                                        //       (terminated)
		.master_burstcount       (),                                        //       (terminated)
		.control_write_base      (26'b00000000000000000000000000),          //       (terminated)
		.control_write_length    (26'b00000000000000000000000000),          //       (terminated)
		.user_write_buffer       (1'b0),                                    //       (terminated)
		.user_buffer_input_data  (32'b00000000000000000000000000000000),    //       (terminated)
		.user_buffer_full        ()                                         //       (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (26),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (26),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) write_master_avalon_master_translator (
		.clk                      (clk_clk),                                                                       //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                //                     reset.reset
		.uav_address              (write_master_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (write_master_avalon_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (write_master_avalon_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (write_master_avalon_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (write_master_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (write_master_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (write_master_avalon_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (write_master_avalon_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (write_master_avalon_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (write_master_avalon_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (write_master_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (write_master_avalon_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (write_master_avalon_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (write_master_avalon_master_byteenable),                                         //                          .byteenable
		.av_write                 (write_master_avalon_master_write),                                              //                          .write
		.av_writedata             (write_master_avalon_master_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                          //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                          //               (terminated)
		.av_begintransfer         (1'b0),                                                                          //               (terminated)
		.av_chipselect            (1'b0),                                                                          //               (terminated)
		.av_read                  (1'b0),                                                                          //               (terminated)
		.av_readdata              (),                                                                              //               (terminated)
		.av_readdatavalid         (),                                                                              //               (terminated)
		.av_lock                  (1'b0),                                                                          //               (terminated)
		.av_debugaccess           (1'b0),                                                                          //               (terminated)
		.uav_clken                (),                                                                              //               (terminated)
		.av_clken                 (1'b1),                                                                          //               (terminated)
		.uav_response             (2'b00),                                                                         //               (terminated)
		.av_response              (),                                                                              //               (terminated)
		.uav_writeresponserequest (),                                                                              //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                          //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                          //               (terminated)
		.av_writeresponsevalid    ()                                                                               //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (26),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (26),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) read_master_avalon_master_translator (
		.clk                      (clk_clk),                                                                      //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                               //                     reset.reset
		.uav_address              (read_master_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (read_master_avalon_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (read_master_avalon_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (read_master_avalon_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (read_master_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (read_master_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (read_master_avalon_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (read_master_avalon_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (read_master_avalon_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (read_master_avalon_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (read_master_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (read_master_avalon_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (read_master_avalon_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (read_master_avalon_master_byteenable),                                         //                          .byteenable
		.av_read                  (read_master_avalon_master_read),                                               //                          .read
		.av_readdata              (read_master_avalon_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (read_master_avalon_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount            (1'b1),                                                                         //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                         //               (terminated)
		.av_begintransfer         (1'b0),                                                                         //               (terminated)
		.av_chipselect            (1'b0),                                                                         //               (terminated)
		.av_write                 (1'b0),                                                                         //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                         //               (terminated)
		.av_lock                  (1'b0),                                                                         //               (terminated)
		.av_debugaccess           (1'b0),                                                                         //               (terminated)
		.uav_clken                (),                                                                             //               (terminated)
		.av_clken                 (1'b1),                                                                         //               (terminated)
		.uav_response             (2'b00),                                                                        //               (terminated)
		.av_response              (),                                                                             //               (terminated)
		.uav_writeresponserequest (),                                                                             //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                         //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                         //               (terminated)
		.av_writeresponsevalid    ()                                                                              //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (24),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) new_sdram_controller_0_s1_translator (
		.clk                      (clk_clk),                                                                              //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                       //                    reset.reset
		.uav_address              (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                                     //              (terminated)
		.av_burstcount            (),                                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                                     //              (terminated)
		.av_lock                  (),                                                                                     //              (terminated)
		.av_clken                 (),                                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                                 //              (terminated)
		.av_debugaccess           (),                                                                                     //              (terminated)
		.av_outputenable          (),                                                                                     //              (terminated)
		.uav_response             (),                                                                                     //              (terminated)
		.av_response              (2'b00),                                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                  //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BURST_SIZE_H          (74),
		.PKT_BURST_SIZE_L          (72),
		.PKT_BURST_TYPE_H          (76),
		.PKT_BURST_TYPE_L          (75),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_TRANS_EXCLUSIVE       (67),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (81),
		.PKT_SRC_ID_L              (81),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (82),
		.PKT_THREAD_ID_H           (83),
		.PKT_THREAD_ID_L           (83),
		.PKT_CACHE_H               (90),
		.PKT_CACHE_L               (87),
		.PKT_DATA_SIDEBAND_H       (78),
		.PKT_DATA_SIDEBAND_L       (78),
		.PKT_QOS_H                 (80),
		.PKT_QOS_L                 (80),
		.PKT_ADDR_SIDEBAND_H       (77),
		.PKT_ADDR_SIDEBAND_L       (77),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.ST_DATA_W                 (93),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) write_master_avalon_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                                //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.av_address              (write_master_avalon_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (write_master_avalon_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (write_master_avalon_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (write_master_avalon_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (write_master_avalon_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (write_master_avalon_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (write_master_avalon_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (write_master_avalon_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (write_master_avalon_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (write_master_avalon_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (write_master_avalon_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (write_master_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (write_master_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (write_master_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (write_master_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (write_master_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_src0_valid),                                                              //        rp.valid
		.rp_data                 (rsp_xbar_demux_src0_data),                                                               //          .data
		.rp_channel              (rsp_xbar_demux_src0_channel),                                                            //          .channel
		.rp_startofpacket        (rsp_xbar_demux_src0_startofpacket),                                                      //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_src0_endofpacket),                                                        //          .endofpacket
		.rp_ready                (rsp_xbar_demux_src0_ready),                                                              //          .ready
		.av_response             (),                                                                                       // (terminated)
		.av_writeresponserequest (1'b0),                                                                                   // (terminated)
		.av_writeresponsevalid   ()                                                                                        // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_BEGIN_BURST           (79),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BURST_SIZE_H          (74),
		.PKT_BURST_SIZE_L          (72),
		.PKT_BURST_TYPE_H          (76),
		.PKT_BURST_TYPE_L          (75),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_TRANS_EXCLUSIVE       (67),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (81),
		.PKT_SRC_ID_L              (81),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (82),
		.PKT_THREAD_ID_H           (83),
		.PKT_THREAD_ID_L           (83),
		.PKT_CACHE_H               (90),
		.PKT_CACHE_L               (87),
		.PKT_DATA_SIDEBAND_H       (78),
		.PKT_DATA_SIDEBAND_L       (78),
		.PKT_QOS_H                 (80),
		.PKT_QOS_L                 (80),
		.PKT_ADDR_SIDEBAND_H       (77),
		.PKT_ADDR_SIDEBAND_L       (77),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.ST_DATA_W                 (93),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) read_master_avalon_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                               //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.av_address              (read_master_avalon_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (read_master_avalon_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (read_master_avalon_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (read_master_avalon_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (read_master_avalon_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (read_master_avalon_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (read_master_avalon_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (read_master_avalon_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (read_master_avalon_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (read_master_avalon_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (read_master_avalon_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (read_master_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (read_master_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (read_master_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (read_master_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (read_master_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_src1_valid),                                                             //        rp.valid
		.rp_data                 (rsp_xbar_demux_src1_data),                                                              //          .data
		.rp_channel              (rsp_xbar_demux_src1_channel),                                                           //          .channel
		.rp_startofpacket        (rsp_xbar_demux_src1_startofpacket),                                                     //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_src1_endofpacket),                                                       //          .endofpacket
		.rp_ready                (rsp_xbar_demux_src1_ready),                                                             //          .ready
		.av_response             (),                                                                                      // (terminated)
		.av_writeresponserequest (1'b0),                                                                                  // (terminated)
		.av_writeresponsevalid   ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (79),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (81),
		.PKT_SRC_ID_L              (81),
		.PKT_DEST_ID_H             (82),
		.PKT_DEST_ID_L             (82),
		.PKT_BURSTWRAP_H           (71),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (86),
		.PKT_PROTECTION_L          (84),
		.PKT_RESPONSE_STATUS_H     (92),
		.PKT_RESPONSE_STATUS_L     (91),
		.PKT_BURST_SIZE_H          (74),
		.PKT_BURST_SIZE_L          (72),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (93),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                         //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                         //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                          //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                       //                .channel
		.rf_sink_ready           (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (94),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                           // (terminated)
		.csr_readdata      (),                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                           // (terminated)
		.almost_full_data  (),                                                                                               // (terminated)
		.almost_empty_data (),                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                           // (terminated)
		.out_empty         (),                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                           // (terminated)
		.out_error         (),                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                           // (terminated)
		.out_channel       ()                                                                                                // (terminated)
	);

	amm_master_qsys_addr_router addr_router (
		.sink_ready         (write_master_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (write_master_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (write_master_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (write_master_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (write_master_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                  //       src.ready
		.src_valid          (addr_router_src_valid),                                                                  //          .valid
		.src_data           (addr_router_src_data),                                                                   //          .data
		.src_channel        (addr_router_src_channel),                                                                //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                             //          .endofpacket
	);

	amm_master_qsys_addr_router addr_router_001 (
		.sink_ready         (read_master_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (read_master_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (read_master_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (read_master_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (read_master_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                             //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                             //          .valid
		.src_data           (addr_router_001_src_data),                                                              //          .data
		.src_channel        (addr_router_001_src_channel),                                                           //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                        //          .endofpacket
	);

	amm_master_qsys_id_router id_router (
		.sink_ready         (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_src_valid),                                                                  //          .valid
		.src_data           (id_router_src_data),                                                                   //          .data
		.src_channel        (id_router_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                             //          .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	amm_master_qsys_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket)    //          .endofpacket
	);

	amm_master_qsys_cmd_xbar_demux cmd_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	amm_master_qsys_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	amm_master_qsys_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

endmodule
