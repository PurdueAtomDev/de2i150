// amm_master_qsys_tb.v

// Generated using ACDS version 13.0sp1 232 at 2014.11.03.12:21:06

`timescale 1 ps / 1 ps
module amm_master_qsys_tb (
	);

	wire    amm_master_qsys_inst_clk_bfm_clk_clk;       // amm_master_qsys_inst_clk_bfm:clk -> [amm_master_qsys_inst:clk_clk, amm_master_qsys_inst_reset_bfm:clk]
	wire    amm_master_qsys_inst_reset_bfm_reset_reset; // amm_master_qsys_inst_reset_bfm:reset -> amm_master_qsys_inst:reset_reset_n

	amm_master_qsys amm_master_qsys_inst (
		.clk_clk                             (amm_master_qsys_inst_clk_bfm_clk_clk),       //                         clk.clk
		.reset_reset_n                       (amm_master_qsys_inst_reset_bfm_reset_reset), //                       reset.reset_n
		.new_sdram_controller_0_wire_addr    (),                                           // new_sdram_controller_0_wire.addr
		.new_sdram_controller_0_wire_ba      (),                                           //                            .ba
		.new_sdram_controller_0_wire_cas_n   (),                                           //                            .cas_n
		.new_sdram_controller_0_wire_cke     (),                                           //                            .cke
		.new_sdram_controller_0_wire_cs_n    (),                                           //                            .cs_n
		.new_sdram_controller_0_wire_dq      (),                                           //                            .dq
		.new_sdram_controller_0_wire_dqm     (),                                           //                            .dqm
		.new_sdram_controller_0_wire_ras_n   (),                                           //                            .ras_n
		.new_sdram_controller_0_wire_we_n    (),                                           //                            .we_n
		.write_master_control_fixed_location (),                                           //        write_master_control.fixed_location
		.write_master_control_write_base     (),                                           //                            .write_base
		.write_master_control_write_length   (),                                           //                            .write_length
		.write_master_control_go             (),                                           //                            .go
		.write_master_control_done           (),                                           //                            .done
		.write_master_user_write_buffer      (),                                           //           write_master_user.write_buffer
		.write_master_user_buffer_input_data (),                                           //                            .buffer_input_data
		.write_master_user_buffer_full       (),                                           //                            .buffer_full
		.read_master_control_fixed_location  (),                                           //         read_master_control.fixed_location
		.read_master_control_read_base       (),                                           //                            .read_base
		.read_master_control_read_length     (),                                           //                            .read_length
		.read_master_control_go              (),                                           //                            .go
		.read_master_control_done            (),                                           //                            .done
		.read_master_control_early_done      (),                                           //                            .early_done
		.read_master_user_read_buffer        (),                                           //            read_master_user.read_buffer
		.read_master_user_buffer_output_data (),                                           //                            .buffer_output_data
		.read_master_user_data_available     ()                                            //                            .data_available
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) amm_master_qsys_inst_clk_bfm (
		.clk (amm_master_qsys_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) amm_master_qsys_inst_reset_bfm (
		.reset (amm_master_qsys_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (amm_master_qsys_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
