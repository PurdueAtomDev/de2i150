// amm_master_qsys_custom_with_bfm_tb.v

// Generated using ACDS version 13.0sp1 232 at 2015.04.20.18:00:05

`timescale 1 ps / 1 ps
module amm_master_qsys_custom_with_bfm_tb (
	);

	wire         amm_master_qsys_custom_with_bfm_inst_clk_bfm_clk_clk;                                // amm_master_qsys_custom_with_bfm_inst_clk_bfm:clk -> [amm_master_qsys_custom_with_bfm_inst:clk_clk, amm_master_qsys_custom_with_bfm_inst_custom_module_conduit_bfm:clk, amm_master_qsys_custom_with_bfm_inst_reset_bfm:clk]
	wire         amm_master_qsys_custom_with_bfm_inst_reset_bfm_reset_reset;                          // amm_master_qsys_custom_with_bfm_inst_reset_bfm:reset -> [amm_master_qsys_custom_with_bfm_inst:reset_reset_n, amm_master_qsys_custom_with_bfm_inst_custom_module_conduit_bfm:reset]
	wire         amm_master_qsys_custom_with_bfm_inst_custom_module_conduit_bfm_conduit_add_data_sel; // amm_master_qsys_custom_with_bfm_inst_custom_module_conduit_bfm:sig_add_data_sel -> amm_master_qsys_custom_with_bfm_inst:custom_module_conduit_add_data_sel
	wire         amm_master_qsys_custom_with_bfm_inst_custom_module_conduit_bfm_conduit_n_action;     // amm_master_qsys_custom_with_bfm_inst_custom_module_conduit_bfm:sig_n_action -> amm_master_qsys_custom_with_bfm_inst:custom_module_conduit_n_action
	wire  [25:0] amm_master_qsys_custom_with_bfm_inst_custom_module_conduit_display_data;             // amm_master_qsys_custom_with_bfm_inst:custom_module_conduit_display_data -> amm_master_qsys_custom_with_bfm_inst_custom_module_conduit_bfm:sig_display_data
	wire         amm_master_qsys_custom_with_bfm_inst_custom_module_conduit_bfm_conduit_rdwr_cntl;    // amm_master_qsys_custom_with_bfm_inst_custom_module_conduit_bfm:sig_rdwr_cntl -> amm_master_qsys_custom_with_bfm_inst:custom_module_conduit_rdwr_cntl
	wire  [25:0] amm_master_qsys_custom_with_bfm_inst_custom_module_conduit_bfm_conduit_rdwr_address; // amm_master_qsys_custom_with_bfm_inst_custom_module_conduit_bfm:sig_rdwr_address -> amm_master_qsys_custom_with_bfm_inst:custom_module_conduit_rdwr_address

	amm_master_qsys_custom_with_bfm amm_master_qsys_custom_with_bfm_inst (
		.clk_clk                            (amm_master_qsys_custom_with_bfm_inst_clk_bfm_clk_clk),                                //                   clk.clk
		.reset_reset_n                      (amm_master_qsys_custom_with_bfm_inst_reset_bfm_reset_reset),                          //                 reset.reset_n
		.custom_module_conduit_rdwr_cntl    (amm_master_qsys_custom_with_bfm_inst_custom_module_conduit_bfm_conduit_rdwr_cntl),    // custom_module_conduit.rdwr_cntl
		.custom_module_conduit_add_data_sel (amm_master_qsys_custom_with_bfm_inst_custom_module_conduit_bfm_conduit_add_data_sel), //                      .add_data_sel
		.custom_module_conduit_rdwr_address (amm_master_qsys_custom_with_bfm_inst_custom_module_conduit_bfm_conduit_rdwr_address), //                      .rdwr_address
		.custom_module_conduit_n_action     (amm_master_qsys_custom_with_bfm_inst_custom_module_conduit_bfm_conduit_n_action),     //                      .n_action
		.custom_module_conduit_display_data (amm_master_qsys_custom_with_bfm_inst_custom_module_conduit_display_data)              //                      .display_data
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) amm_master_qsys_custom_with_bfm_inst_clk_bfm (
		.clk (amm_master_qsys_custom_with_bfm_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) amm_master_qsys_custom_with_bfm_inst_reset_bfm (
		.reset (amm_master_qsys_custom_with_bfm_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (amm_master_qsys_custom_with_bfm_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm amm_master_qsys_custom_with_bfm_inst_custom_module_conduit_bfm (
		.clk              (amm_master_qsys_custom_with_bfm_inst_clk_bfm_clk_clk),                                //     clk.clk
		.reset            (~amm_master_qsys_custom_with_bfm_inst_reset_bfm_reset_reset),                         //   reset.reset
		.sig_rdwr_cntl    (amm_master_qsys_custom_with_bfm_inst_custom_module_conduit_bfm_conduit_rdwr_cntl),    // conduit.rdwr_cntl
		.sig_add_data_sel (amm_master_qsys_custom_with_bfm_inst_custom_module_conduit_bfm_conduit_add_data_sel), //        .add_data_sel
		.sig_rdwr_address (amm_master_qsys_custom_with_bfm_inst_custom_module_conduit_bfm_conduit_rdwr_address), //        .rdwr_address
		.sig_n_action     (amm_master_qsys_custom_with_bfm_inst_custom_module_conduit_bfm_conduit_n_action),     //        .n_action
		.sig_display_data (amm_master_qsys_custom_with_bfm_inst_custom_module_conduit_display_data)              //        .display_data
	);

endmodule
