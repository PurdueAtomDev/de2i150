// amm_master_qsys_with_pcie.v

// Generated using ACDS version 13.0sp1 232 at 2015.03.31.16:42:38

`timescale 1 ps / 1 ps
module amm_master_qsys_with_pcie (
		input  wire        clk_clk,                                    //                        clk.clk
		input  wire        reset_reset_n,                              //                      reset.reset_n
		input  wire [3:0]  pcie_ip_reconfig_togxb_data,                //     pcie_ip_reconfig_togxb.data
		input  wire        pcie_ip_refclk_export,                      //             pcie_ip_refclk.export
		input  wire [39:0] pcie_ip_test_in_test_in,                    //            pcie_ip_test_in.test_in
		input  wire        pcie_ip_pcie_rstn_export,                   //          pcie_ip_pcie_rstn.export
		output wire        pcie_ip_clocks_sim_clk250_export,           //         pcie_ip_clocks_sim.clk250_export
		output wire        pcie_ip_clocks_sim_clk500_export,           //                           .clk500_export
		output wire        pcie_ip_clocks_sim_clk125_export,           //                           .clk125_export
		input  wire        pcie_ip_reconfig_busy_busy_altgxb_reconfig, //      pcie_ip_reconfig_busy.busy_altgxb_reconfig
		input  wire        pcie_ip_pipe_ext_pipe_mode,                 //           pcie_ip_pipe_ext.pipe_mode
		input  wire        pcie_ip_pipe_ext_phystatus_ext,             //                           .phystatus_ext
		output wire        pcie_ip_pipe_ext_rate_ext,                  //                           .rate_ext
		output wire [1:0]  pcie_ip_pipe_ext_powerdown_ext,             //                           .powerdown_ext
		output wire        pcie_ip_pipe_ext_txdetectrx_ext,            //                           .txdetectrx_ext
		input  wire        pcie_ip_pipe_ext_rxelecidle0_ext,           //                           .rxelecidle0_ext
		input  wire [7:0]  pcie_ip_pipe_ext_rxdata0_ext,               //                           .rxdata0_ext
		input  wire [2:0]  pcie_ip_pipe_ext_rxstatus0_ext,             //                           .rxstatus0_ext
		input  wire        pcie_ip_pipe_ext_rxvalid0_ext,              //                           .rxvalid0_ext
		input  wire        pcie_ip_pipe_ext_rxdatak0_ext,              //                           .rxdatak0_ext
		output wire [7:0]  pcie_ip_pipe_ext_txdata0_ext,               //                           .txdata0_ext
		output wire        pcie_ip_pipe_ext_txdatak0_ext,              //                           .txdatak0_ext
		output wire        pcie_ip_pipe_ext_rxpolarity0_ext,           //                           .rxpolarity0_ext
		output wire        pcie_ip_pipe_ext_txcompl0_ext,              //                           .txcompl0_ext
		output wire        pcie_ip_pipe_ext_txelecidle0_ext,           //                           .txelecidle0_ext
		input  wire        pcie_ip_rx_in_rx_datain_0,                  //              pcie_ip_rx_in.rx_datain_0
		output wire        pcie_ip_tx_out_tx_dataout_0,                //             pcie_ip_tx_out.tx_dataout_0
		output wire [4:0]  pcie_ip_reconfig_fromgxb_0_data,            // pcie_ip_reconfig_fromgxb_0.data
		output wire [11:0] sdram_addr,                                 //                      sdram.addr
		output wire [1:0]  sdram_ba,                                   //                           .ba
		output wire        sdram_cas_n,                                //                           .cas_n
		output wire        sdram_cke,                                  //                           .cke
		output wire        sdram_cs_n,                                 //                           .cs_n
		inout  wire [31:0] sdram_dq,                                   //                           .dq
		output wire [3:0]  sdram_dqm,                                  //                           .dqm
		output wire        sdram_ras_n,                                //                           .ras_n
		output wire        sdram_we_n,                                 //                           .we_n
		output wire        altpll_sdram_clk,                           //               altpll_sdram.clk
		input  wire        pcie_ip_powerdown_pll_powerdown,            //          pcie_ip_powerdown.pll_powerdown
		input  wire        pcie_ip_powerdown_gxb_powerdown,            //                           .gxb_powerdown
		input  wire        custom_module_conduit_rdwr_cntl,            //      custom_module_conduit.rdwr_cntl
		input  wire        custom_module_conduit_n_action,             //                           .n_action
		input  wire        custom_module_conduit_add_data_sel,         //                           .add_data_sel
		input  wire [27:0] custom_module_conduit_rdwr_address          //                           .rdwr_address
	);

	wire          pcie_ip_pcie_core_clk_clk;                                                                              // pcie_ip:pcie_core_clk_clk -> [addr_router:clk, addr_router_001:clk, addr_router_002:clk, addr_router_003:clk, addr_router_004:clk, addr_router_005:clk, burst_adapter:clk, burst_adapter_001:clk, burst_adapter_002:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_demux_002:clk, cmd_xbar_demux_003:clk, cmd_xbar_demux_004:clk, cmd_xbar_demux_005:clk, cmd_xbar_mux_002:clk, crosser:in_clk, crosser_001:out_clk, crosser_002:in_clk, crosser_003:in_clk, crosser_004:out_clk, crosser_005:out_clk, id_router:clk, id_router_001:clk, id_router_002:clk, irq_mapper:clk, limiter:clk, limiter_001:clk, pcie_ip:fixedclk_clk, pcie_ip_bar1_0_translator:clk, pcie_ip_bar1_0_translator_avalon_universal_master_0_agent:clk, pcie_ip_bar2_translator:clk, pcie_ip_bar2_translator_avalon_universal_master_0_agent:clk, pcie_ip_cra_translator:clk, pcie_ip_cra_translator_avalon_universal_slave_0_agent:clk, pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pcie_ip_txs_translator:clk, pcie_ip_txs_translator_avalon_universal_slave_0_agent:clk, pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_mux:clk, rsp_xbar_mux_003:clk, rsp_xbar_mux_004:clk, rst_controller:clk, rst_controller_003:clk, sgdma:clk, sgdma_csr_translator:clk, sgdma_csr_translator_avalon_universal_slave_0_agent:clk, sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sgdma_descriptor_read_translator:clk, sgdma_descriptor_read_translator_avalon_universal_master_0_agent:clk, sgdma_descriptor_write_translator:clk, sgdma_descriptor_write_translator_avalon_universal_master_0_agent:clk, sgdma_m_read_translator:clk, sgdma_m_read_translator_avalon_universal_master_0_agent:clk, sgdma_m_write_translator:clk, sgdma_m_write_translator_avalon_universal_master_0_agent:clk, width_adapter:clk, width_adapter_001:clk, width_adapter_002:clk, width_adapter_003:clk, width_adapter_004:clk, width_adapter_005:clk, width_adapter_006:clk, width_adapter_007:clk, width_adapter_008:clk, width_adapter_009:clk]
	wire          altpll_qsys_c3_clk;                                                                                     // altpll_qsys:c3 -> [pcie_ip:cal_blk_clk_clk, pcie_ip:reconfig_gxbclk_clk]
	wire    [6:0] pcie_ip_bar2_burstcount;                                                                                // pcie_ip:bar2_burstcount -> pcie_ip_bar2_translator:av_burstcount
	wire          pcie_ip_bar2_waitrequest;                                                                               // pcie_ip_bar2_translator:av_waitrequest -> pcie_ip:bar2_waitrequest
	wire   [63:0] pcie_ip_bar2_writedata;                                                                                 // pcie_ip:bar2_writedata -> pcie_ip_bar2_translator:av_writedata
	wire   [31:0] pcie_ip_bar2_address;                                                                                   // pcie_ip:bar2_address -> pcie_ip_bar2_translator:av_address
	wire          pcie_ip_bar2_write;                                                                                     // pcie_ip:bar2_write -> pcie_ip_bar2_translator:av_write
	wire          pcie_ip_bar2_read;                                                                                      // pcie_ip:bar2_read -> pcie_ip_bar2_translator:av_read
	wire   [63:0] pcie_ip_bar2_readdata;                                                                                  // pcie_ip_bar2_translator:av_readdata -> pcie_ip:bar2_readdata
	wire    [7:0] pcie_ip_bar2_byteenable;                                                                                // pcie_ip:bar2_byteenable -> pcie_ip_bar2_translator:av_byteenable
	wire          pcie_ip_bar2_readdatavalid;                                                                             // pcie_ip_bar2_translator:av_readdatavalid -> pcie_ip:bar2_readdatavalid
	wire   [31:0] sgdma_csr_translator_avalon_anti_slave_0_writedata;                                                     // sgdma_csr_translator:av_writedata -> sgdma:csr_writedata
	wire    [3:0] sgdma_csr_translator_avalon_anti_slave_0_address;                                                       // sgdma_csr_translator:av_address -> sgdma:csr_address
	wire          sgdma_csr_translator_avalon_anti_slave_0_chipselect;                                                    // sgdma_csr_translator:av_chipselect -> sgdma:csr_chipselect
	wire          sgdma_csr_translator_avalon_anti_slave_0_write;                                                         // sgdma_csr_translator:av_write -> sgdma:csr_write
	wire          sgdma_csr_translator_avalon_anti_slave_0_read;                                                          // sgdma_csr_translator:av_read -> sgdma:csr_read
	wire   [31:0] sgdma_csr_translator_avalon_anti_slave_0_readdata;                                                      // sgdma:csr_readdata -> sgdma_csr_translator:av_readdata
	wire          pcie_ip_cra_translator_avalon_anti_slave_0_waitrequest;                                                 // pcie_ip:cra_waitrequest -> pcie_ip_cra_translator:av_waitrequest
	wire   [31:0] pcie_ip_cra_translator_avalon_anti_slave_0_writedata;                                                   // pcie_ip_cra_translator:av_writedata -> pcie_ip:cra_writedata
	wire   [11:0] pcie_ip_cra_translator_avalon_anti_slave_0_address;                                                     // pcie_ip_cra_translator:av_address -> pcie_ip:cra_address
	wire          pcie_ip_cra_translator_avalon_anti_slave_0_chipselect;                                                  // pcie_ip_cra_translator:av_chipselect -> pcie_ip:cra_chipselect
	wire          pcie_ip_cra_translator_avalon_anti_slave_0_write;                                                       // pcie_ip_cra_translator:av_write -> pcie_ip:cra_write
	wire          pcie_ip_cra_translator_avalon_anti_slave_0_read;                                                        // pcie_ip_cra_translator:av_read -> pcie_ip:cra_read
	wire   [31:0] pcie_ip_cra_translator_avalon_anti_slave_0_readdata;                                                    // pcie_ip:cra_readdata -> pcie_ip_cra_translator:av_readdata
	wire    [3:0] pcie_ip_cra_translator_avalon_anti_slave_0_byteenable;                                                  // pcie_ip_cra_translator:av_byteenable -> pcie_ip:cra_byteenable
	wire          sgdma_descriptor_read_waitrequest;                                                                      // sgdma_descriptor_read_translator:av_waitrequest -> sgdma:descriptor_read_waitrequest
	wire   [31:0] sgdma_descriptor_read_address;                                                                          // sgdma:descriptor_read_address -> sgdma_descriptor_read_translator:av_address
	wire          sgdma_descriptor_read_read;                                                                             // sgdma:descriptor_read_read -> sgdma_descriptor_read_translator:av_read
	wire   [31:0] sgdma_descriptor_read_readdata;                                                                         // sgdma_descriptor_read_translator:av_readdata -> sgdma:descriptor_read_readdata
	wire          sgdma_descriptor_read_readdatavalid;                                                                    // sgdma_descriptor_read_translator:av_readdatavalid -> sgdma:descriptor_read_readdatavalid
	wire          sgdma_descriptor_write_waitrequest;                                                                     // sgdma_descriptor_write_translator:av_waitrequest -> sgdma:descriptor_write_waitrequest
	wire   [31:0] sgdma_descriptor_write_writedata;                                                                       // sgdma:descriptor_write_writedata -> sgdma_descriptor_write_translator:av_writedata
	wire   [31:0] sgdma_descriptor_write_address;                                                                         // sgdma:descriptor_write_address -> sgdma_descriptor_write_translator:av_address
	wire          sgdma_descriptor_write_write;                                                                           // sgdma:descriptor_write_write -> sgdma_descriptor_write_translator:av_write
	wire    [3:0] sgdma_m_read_burstcount;                                                                                // sgdma:m_read_burstcount -> sgdma_m_read_translator:av_burstcount
	wire          sgdma_m_read_waitrequest;                                                                               // sgdma_m_read_translator:av_waitrequest -> sgdma:m_read_waitrequest
	wire   [31:0] sgdma_m_read_address;                                                                                   // sgdma:m_read_address -> sgdma_m_read_translator:av_address
	wire          sgdma_m_read_read;                                                                                      // sgdma:m_read_read -> sgdma_m_read_translator:av_read
	wire   [63:0] sgdma_m_read_readdata;                                                                                  // sgdma_m_read_translator:av_readdata -> sgdma:m_read_readdata
	wire          sgdma_m_read_readdatavalid;                                                                             // sgdma_m_read_translator:av_readdatavalid -> sgdma:m_read_readdatavalid
	wire    [7:0] sgdma_m_write_burstcount;                                                                               // sgdma:m_write_burstcount -> sgdma_m_write_translator:av_burstcount
	wire          sgdma_m_write_waitrequest;                                                                              // sgdma_m_write_translator:av_waitrequest -> sgdma:m_write_waitrequest
	wire   [63:0] sgdma_m_write_writedata;                                                                                // sgdma:m_write_writedata -> sgdma_m_write_translator:av_writedata
	wire   [31:0] sgdma_m_write_address;                                                                                  // sgdma:m_write_address -> sgdma_m_write_translator:av_address
	wire          sgdma_m_write_write;                                                                                    // sgdma:m_write_write -> sgdma_m_write_translator:av_write
	wire    [7:0] sgdma_m_write_byteenable;                                                                               // sgdma:m_write_byteenable -> sgdma_m_write_translator:av_byteenable
	wire          pcie_ip_txs_translator_avalon_anti_slave_0_waitrequest;                                                 // pcie_ip:txs_waitrequest -> pcie_ip_txs_translator:av_waitrequest
	wire    [6:0] pcie_ip_txs_translator_avalon_anti_slave_0_burstcount;                                                  // pcie_ip_txs_translator:av_burstcount -> pcie_ip:txs_burstcount
	wire   [63:0] pcie_ip_txs_translator_avalon_anti_slave_0_writedata;                                                   // pcie_ip_txs_translator:av_writedata -> pcie_ip:txs_writedata
	wire   [30:0] pcie_ip_txs_translator_avalon_anti_slave_0_address;                                                     // pcie_ip_txs_translator:av_address -> pcie_ip:txs_address
	wire          pcie_ip_txs_translator_avalon_anti_slave_0_chipselect;                                                  // pcie_ip_txs_translator:av_chipselect -> pcie_ip:txs_chipselect
	wire          pcie_ip_txs_translator_avalon_anti_slave_0_write;                                                       // pcie_ip_txs_translator:av_write -> pcie_ip:txs_write
	wire          pcie_ip_txs_translator_avalon_anti_slave_0_read;                                                        // pcie_ip_txs_translator:av_read -> pcie_ip:txs_read
	wire   [63:0] pcie_ip_txs_translator_avalon_anti_slave_0_readdata;                                                    // pcie_ip:txs_readdata -> pcie_ip_txs_translator:av_readdata
	wire          pcie_ip_txs_translator_avalon_anti_slave_0_readdatavalid;                                               // pcie_ip:txs_readdatavalid -> pcie_ip_txs_translator:av_readdatavalid
	wire    [7:0] pcie_ip_txs_translator_avalon_anti_slave_0_byteenable;                                                  // pcie_ip_txs_translator:av_byteenable -> pcie_ip:txs_byteenable
	wire          sdram_s1_translator_avalon_anti_slave_0_waitrequest;                                                    // sdram:za_waitrequest -> sdram_s1_translator:av_waitrequest
	wire   [31:0] sdram_s1_translator_avalon_anti_slave_0_writedata;                                                      // sdram_s1_translator:av_writedata -> sdram:az_data
	wire   [23:0] sdram_s1_translator_avalon_anti_slave_0_address;                                                        // sdram_s1_translator:av_address -> sdram:az_addr
	wire          sdram_s1_translator_avalon_anti_slave_0_chipselect;                                                     // sdram_s1_translator:av_chipselect -> sdram:az_cs
	wire          sdram_s1_translator_avalon_anti_slave_0_write;                                                          // sdram_s1_translator:av_write -> sdram:az_wr_n
	wire          sdram_s1_translator_avalon_anti_slave_0_read;                                                           // sdram_s1_translator:av_read -> sdram:az_rd_n
	wire   [31:0] sdram_s1_translator_avalon_anti_slave_0_readdata;                                                       // sdram:za_data -> sdram_s1_translator:av_readdata
	wire          sdram_s1_translator_avalon_anti_slave_0_readdatavalid;                                                  // sdram:za_valid -> sdram_s1_translator:av_readdatavalid
	wire    [3:0] sdram_s1_translator_avalon_anti_slave_0_byteenable;                                                     // sdram_s1_translator:av_byteenable -> sdram:az_be_n
	wire    [6:0] pcie_ip_bar1_0_burstcount;                                                                              // pcie_ip:bar1_0_burstcount -> pcie_ip_bar1_0_translator:av_burstcount
	wire          pcie_ip_bar1_0_waitrequest;                                                                             // pcie_ip_bar1_0_translator:av_waitrequest -> pcie_ip:bar1_0_waitrequest
	wire   [63:0] pcie_ip_bar1_0_writedata;                                                                               // pcie_ip:bar1_0_writedata -> pcie_ip_bar1_0_translator:av_writedata
	wire   [31:0] pcie_ip_bar1_0_address;                                                                                 // pcie_ip:bar1_0_address -> pcie_ip_bar1_0_translator:av_address
	wire          pcie_ip_bar1_0_write;                                                                                   // pcie_ip:bar1_0_write -> pcie_ip_bar1_0_translator:av_write
	wire          pcie_ip_bar1_0_read;                                                                                    // pcie_ip:bar1_0_read -> pcie_ip_bar1_0_translator:av_read
	wire   [63:0] pcie_ip_bar1_0_readdata;                                                                                // pcie_ip_bar1_0_translator:av_readdata -> pcie_ip:bar1_0_readdata
	wire    [7:0] pcie_ip_bar1_0_byteenable;                                                                              // pcie_ip:bar1_0_byteenable -> pcie_ip_bar1_0_translator:av_byteenable
	wire          pcie_ip_bar1_0_readdatavalid;                                                                           // pcie_ip_bar1_0_translator:av_readdatavalid -> pcie_ip:bar1_0_readdatavalid
	wire   [31:0] custom_slave_block_0_avalon_slave_translator_avalon_anti_slave_0_writedata;                             // custom_slave_block_0_avalon_slave_translator:av_writedata -> custom_slave_block_0:slave_writedata
	wire    [4:0] custom_slave_block_0_avalon_slave_translator_avalon_anti_slave_0_address;                               // custom_slave_block_0_avalon_slave_translator:av_address -> custom_slave_block_0:slave_address
	wire          custom_slave_block_0_avalon_slave_translator_avalon_anti_slave_0_chipselect;                            // custom_slave_block_0_avalon_slave_translator:av_chipselect -> custom_slave_block_0:slave_chipselect
	wire          custom_slave_block_0_avalon_slave_translator_avalon_anti_slave_0_write;                                 // custom_slave_block_0_avalon_slave_translator:av_write -> custom_slave_block_0:slave_write
	wire          custom_slave_block_0_avalon_slave_translator_avalon_anti_slave_0_read;                                  // custom_slave_block_0_avalon_slave_translator:av_read -> custom_slave_block_0:slave_read
	wire   [31:0] custom_slave_block_0_avalon_slave_translator_avalon_anti_slave_0_readdata;                              // custom_slave_block_0:slave_readdata -> custom_slave_block_0_avalon_slave_translator:av_readdata
	wire          pcie_ip_bar2_translator_avalon_universal_master_0_waitrequest;                                          // pcie_ip_bar2_translator_avalon_universal_master_0_agent:av_waitrequest -> pcie_ip_bar2_translator:uav_waitrequest
	wire    [9:0] pcie_ip_bar2_translator_avalon_universal_master_0_burstcount;                                           // pcie_ip_bar2_translator:uav_burstcount -> pcie_ip_bar2_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [63:0] pcie_ip_bar2_translator_avalon_universal_master_0_writedata;                                            // pcie_ip_bar2_translator:uav_writedata -> pcie_ip_bar2_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] pcie_ip_bar2_translator_avalon_universal_master_0_address;                                              // pcie_ip_bar2_translator:uav_address -> pcie_ip_bar2_translator_avalon_universal_master_0_agent:av_address
	wire          pcie_ip_bar2_translator_avalon_universal_master_0_lock;                                                 // pcie_ip_bar2_translator:uav_lock -> pcie_ip_bar2_translator_avalon_universal_master_0_agent:av_lock
	wire          pcie_ip_bar2_translator_avalon_universal_master_0_write;                                                // pcie_ip_bar2_translator:uav_write -> pcie_ip_bar2_translator_avalon_universal_master_0_agent:av_write
	wire          pcie_ip_bar2_translator_avalon_universal_master_0_read;                                                 // pcie_ip_bar2_translator:uav_read -> pcie_ip_bar2_translator_avalon_universal_master_0_agent:av_read
	wire   [63:0] pcie_ip_bar2_translator_avalon_universal_master_0_readdata;                                             // pcie_ip_bar2_translator_avalon_universal_master_0_agent:av_readdata -> pcie_ip_bar2_translator:uav_readdata
	wire          pcie_ip_bar2_translator_avalon_universal_master_0_debugaccess;                                          // pcie_ip_bar2_translator:uav_debugaccess -> pcie_ip_bar2_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [7:0] pcie_ip_bar2_translator_avalon_universal_master_0_byteenable;                                           // pcie_ip_bar2_translator:uav_byteenable -> pcie_ip_bar2_translator_avalon_universal_master_0_agent:av_byteenable
	wire          pcie_ip_bar2_translator_avalon_universal_master_0_readdatavalid;                                        // pcie_ip_bar2_translator_avalon_universal_master_0_agent:av_readdatavalid -> pcie_ip_bar2_translator:uav_readdatavalid
	wire          sgdma_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // sgdma_csr_translator:uav_waitrequest -> sgdma_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sgdma_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // sgdma_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> sgdma_csr_translator:uav_burstcount
	wire   [31:0] sgdma_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // sgdma_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> sgdma_csr_translator:uav_writedata
	wire   [31:0] sgdma_csr_translator_avalon_universal_slave_0_agent_m0_address;                                         // sgdma_csr_translator_avalon_universal_slave_0_agent:m0_address -> sgdma_csr_translator:uav_address
	wire          sgdma_csr_translator_avalon_universal_slave_0_agent_m0_write;                                           // sgdma_csr_translator_avalon_universal_slave_0_agent:m0_write -> sgdma_csr_translator:uav_write
	wire          sgdma_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                            // sgdma_csr_translator_avalon_universal_slave_0_agent:m0_lock -> sgdma_csr_translator:uav_lock
	wire          sgdma_csr_translator_avalon_universal_slave_0_agent_m0_read;                                            // sgdma_csr_translator_avalon_universal_slave_0_agent:m0_read -> sgdma_csr_translator:uav_read
	wire   [31:0] sgdma_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // sgdma_csr_translator:uav_readdata -> sgdma_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sgdma_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // sgdma_csr_translator:uav_readdatavalid -> sgdma_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sgdma_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // sgdma_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sgdma_csr_translator:uav_debugaccess
	wire    [3:0] sgdma_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // sgdma_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> sgdma_csr_translator:uav_byteenable
	wire          sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // sgdma_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // sgdma_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // sgdma_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [106:0] sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // sgdma_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sgdma_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sgdma_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sgdma_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sgdma_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [106:0] sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sgdma_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // sgdma_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sgdma_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // sgdma_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sgdma_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] sgdma_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // sgdma_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sgdma_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sgdma_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // sgdma_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sgdma_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // pcie_ip_cra_translator:uav_waitrequest -> pcie_ip_cra_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // pcie_ip_cra_translator_avalon_universal_slave_0_agent:m0_burstcount -> pcie_ip_cra_translator:uav_burstcount
	wire   [31:0] pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // pcie_ip_cra_translator_avalon_universal_slave_0_agent:m0_writedata -> pcie_ip_cra_translator:uav_writedata
	wire   [31:0] pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_address;                                       // pcie_ip_cra_translator_avalon_universal_slave_0_agent:m0_address -> pcie_ip_cra_translator:uav_address
	wire          pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_write;                                         // pcie_ip_cra_translator_avalon_universal_slave_0_agent:m0_write -> pcie_ip_cra_translator:uav_write
	wire          pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_lock;                                          // pcie_ip_cra_translator_avalon_universal_slave_0_agent:m0_lock -> pcie_ip_cra_translator:uav_lock
	wire          pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_read;                                          // pcie_ip_cra_translator_avalon_universal_slave_0_agent:m0_read -> pcie_ip_cra_translator:uav_read
	wire   [31:0] pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // pcie_ip_cra_translator:uav_readdata -> pcie_ip_cra_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // pcie_ip_cra_translator:uav_readdatavalid -> pcie_ip_cra_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // pcie_ip_cra_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pcie_ip_cra_translator:uav_debugaccess
	wire    [3:0] pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // pcie_ip_cra_translator_avalon_universal_slave_0_agent:m0_byteenable -> pcie_ip_cra_translator:uav_byteenable
	wire          pcie_ip_cra_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // pcie_ip_cra_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pcie_ip_cra_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // pcie_ip_cra_translator_avalon_universal_slave_0_agent:rf_source_valid -> pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pcie_ip_cra_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // pcie_ip_cra_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [106:0] pcie_ip_cra_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // pcie_ip_cra_translator_avalon_universal_slave_0_agent:rf_source_data -> pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pcie_ip_cra_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pcie_ip_cra_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pcie_ip_cra_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pcie_ip_cra_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pcie_ip_cra_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [106:0] pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pcie_ip_cra_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // pcie_ip_cra_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pcie_ip_cra_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // pcie_ip_cra_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pcie_ip_cra_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] pcie_ip_cra_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // pcie_ip_cra_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pcie_ip_cra_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pcie_ip_cra_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // pcie_ip_cra_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pcie_ip_cra_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sgdma_descriptor_read_translator_avalon_universal_master_0_waitrequest;                                 // sgdma_descriptor_read_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_descriptor_read_translator:uav_waitrequest
	wire    [2:0] sgdma_descriptor_read_translator_avalon_universal_master_0_burstcount;                                  // sgdma_descriptor_read_translator:uav_burstcount -> sgdma_descriptor_read_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_descriptor_read_translator_avalon_universal_master_0_writedata;                                   // sgdma_descriptor_read_translator:uav_writedata -> sgdma_descriptor_read_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_descriptor_read_translator_avalon_universal_master_0_address;                                     // sgdma_descriptor_read_translator:uav_address -> sgdma_descriptor_read_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_descriptor_read_translator_avalon_universal_master_0_lock;                                        // sgdma_descriptor_read_translator:uav_lock -> sgdma_descriptor_read_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_descriptor_read_translator_avalon_universal_master_0_write;                                       // sgdma_descriptor_read_translator:uav_write -> sgdma_descriptor_read_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_descriptor_read_translator_avalon_universal_master_0_read;                                        // sgdma_descriptor_read_translator:uav_read -> sgdma_descriptor_read_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_descriptor_read_translator_avalon_universal_master_0_readdata;                                    // sgdma_descriptor_read_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_descriptor_read_translator:uav_readdata
	wire          sgdma_descriptor_read_translator_avalon_universal_master_0_debugaccess;                                 // sgdma_descriptor_read_translator:uav_debugaccess -> sgdma_descriptor_read_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_descriptor_read_translator_avalon_universal_master_0_byteenable;                                  // sgdma_descriptor_read_translator:uav_byteenable -> sgdma_descriptor_read_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_descriptor_read_translator_avalon_universal_master_0_readdatavalid;                               // sgdma_descriptor_read_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_descriptor_read_translator:uav_readdatavalid
	wire          sgdma_descriptor_write_translator_avalon_universal_master_0_waitrequest;                                // sgdma_descriptor_write_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_descriptor_write_translator:uav_waitrequest
	wire    [2:0] sgdma_descriptor_write_translator_avalon_universal_master_0_burstcount;                                 // sgdma_descriptor_write_translator:uav_burstcount -> sgdma_descriptor_write_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_descriptor_write_translator_avalon_universal_master_0_writedata;                                  // sgdma_descriptor_write_translator:uav_writedata -> sgdma_descriptor_write_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_descriptor_write_translator_avalon_universal_master_0_address;                                    // sgdma_descriptor_write_translator:uav_address -> sgdma_descriptor_write_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_descriptor_write_translator_avalon_universal_master_0_lock;                                       // sgdma_descriptor_write_translator:uav_lock -> sgdma_descriptor_write_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_descriptor_write_translator_avalon_universal_master_0_write;                                      // sgdma_descriptor_write_translator:uav_write -> sgdma_descriptor_write_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_descriptor_write_translator_avalon_universal_master_0_read;                                       // sgdma_descriptor_write_translator:uav_read -> sgdma_descriptor_write_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_descriptor_write_translator_avalon_universal_master_0_readdata;                                   // sgdma_descriptor_write_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_descriptor_write_translator:uav_readdata
	wire          sgdma_descriptor_write_translator_avalon_universal_master_0_debugaccess;                                // sgdma_descriptor_write_translator:uav_debugaccess -> sgdma_descriptor_write_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_descriptor_write_translator_avalon_universal_master_0_byteenable;                                 // sgdma_descriptor_write_translator:uav_byteenable -> sgdma_descriptor_write_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_descriptor_write_translator_avalon_universal_master_0_readdatavalid;                              // sgdma_descriptor_write_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_descriptor_write_translator:uav_readdatavalid
	wire          sgdma_m_read_translator_avalon_universal_master_0_waitrequest;                                          // sgdma_m_read_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_m_read_translator:uav_waitrequest
	wire    [6:0] sgdma_m_read_translator_avalon_universal_master_0_burstcount;                                           // sgdma_m_read_translator:uav_burstcount -> sgdma_m_read_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [63:0] sgdma_m_read_translator_avalon_universal_master_0_writedata;                                            // sgdma_m_read_translator:uav_writedata -> sgdma_m_read_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_m_read_translator_avalon_universal_master_0_address;                                              // sgdma_m_read_translator:uav_address -> sgdma_m_read_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_m_read_translator_avalon_universal_master_0_lock;                                                 // sgdma_m_read_translator:uav_lock -> sgdma_m_read_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_m_read_translator_avalon_universal_master_0_write;                                                // sgdma_m_read_translator:uav_write -> sgdma_m_read_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_m_read_translator_avalon_universal_master_0_read;                                                 // sgdma_m_read_translator:uav_read -> sgdma_m_read_translator_avalon_universal_master_0_agent:av_read
	wire   [63:0] sgdma_m_read_translator_avalon_universal_master_0_readdata;                                             // sgdma_m_read_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_m_read_translator:uav_readdata
	wire          sgdma_m_read_translator_avalon_universal_master_0_debugaccess;                                          // sgdma_m_read_translator:uav_debugaccess -> sgdma_m_read_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [7:0] sgdma_m_read_translator_avalon_universal_master_0_byteenable;                                           // sgdma_m_read_translator:uav_byteenable -> sgdma_m_read_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_m_read_translator_avalon_universal_master_0_readdatavalid;                                        // sgdma_m_read_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_m_read_translator:uav_readdatavalid
	wire          sgdma_m_write_translator_avalon_universal_master_0_waitrequest;                                         // sgdma_m_write_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_m_write_translator:uav_waitrequest
	wire   [10:0] sgdma_m_write_translator_avalon_universal_master_0_burstcount;                                          // sgdma_m_write_translator:uav_burstcount -> sgdma_m_write_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [63:0] sgdma_m_write_translator_avalon_universal_master_0_writedata;                                           // sgdma_m_write_translator:uav_writedata -> sgdma_m_write_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_m_write_translator_avalon_universal_master_0_address;                                             // sgdma_m_write_translator:uav_address -> sgdma_m_write_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_m_write_translator_avalon_universal_master_0_lock;                                                // sgdma_m_write_translator:uav_lock -> sgdma_m_write_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_m_write_translator_avalon_universal_master_0_write;                                               // sgdma_m_write_translator:uav_write -> sgdma_m_write_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_m_write_translator_avalon_universal_master_0_read;                                                // sgdma_m_write_translator:uav_read -> sgdma_m_write_translator_avalon_universal_master_0_agent:av_read
	wire   [63:0] sgdma_m_write_translator_avalon_universal_master_0_readdata;                                            // sgdma_m_write_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_m_write_translator:uav_readdata
	wire          sgdma_m_write_translator_avalon_universal_master_0_debugaccess;                                         // sgdma_m_write_translator:uav_debugaccess -> sgdma_m_write_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [7:0] sgdma_m_write_translator_avalon_universal_master_0_byteenable;                                          // sgdma_m_write_translator:uav_byteenable -> sgdma_m_write_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_m_write_translator_avalon_universal_master_0_readdatavalid;                                       // sgdma_m_write_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_m_write_translator:uav_readdatavalid
	wire          pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // pcie_ip_txs_translator:uav_waitrequest -> pcie_ip_txs_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [9:0] pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // pcie_ip_txs_translator_avalon_universal_slave_0_agent:m0_burstcount -> pcie_ip_txs_translator:uav_burstcount
	wire   [63:0] pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // pcie_ip_txs_translator_avalon_universal_slave_0_agent:m0_writedata -> pcie_ip_txs_translator:uav_writedata
	wire   [31:0] pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_address;                                       // pcie_ip_txs_translator_avalon_universal_slave_0_agent:m0_address -> pcie_ip_txs_translator:uav_address
	wire          pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_write;                                         // pcie_ip_txs_translator_avalon_universal_slave_0_agent:m0_write -> pcie_ip_txs_translator:uav_write
	wire          pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_lock;                                          // pcie_ip_txs_translator_avalon_universal_slave_0_agent:m0_lock -> pcie_ip_txs_translator:uav_lock
	wire          pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_read;                                          // pcie_ip_txs_translator_avalon_universal_slave_0_agent:m0_read -> pcie_ip_txs_translator:uav_read
	wire   [63:0] pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // pcie_ip_txs_translator:uav_readdata -> pcie_ip_txs_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // pcie_ip_txs_translator:uav_readdatavalid -> pcie_ip_txs_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // pcie_ip_txs_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pcie_ip_txs_translator:uav_debugaccess
	wire    [7:0] pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // pcie_ip_txs_translator_avalon_universal_slave_0_agent:m0_byteenable -> pcie_ip_txs_translator:uav_byteenable
	wire          pcie_ip_txs_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // pcie_ip_txs_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pcie_ip_txs_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // pcie_ip_txs_translator_avalon_universal_slave_0_agent:rf_source_valid -> pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pcie_ip_txs_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // pcie_ip_txs_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [145:0] pcie_ip_txs_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // pcie_ip_txs_translator_avalon_universal_slave_0_agent:rf_source_data -> pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pcie_ip_txs_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pcie_ip_txs_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pcie_ip_txs_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pcie_ip_txs_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pcie_ip_txs_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [145:0] pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pcie_ip_txs_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // pcie_ip_txs_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pcie_ip_txs_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // pcie_ip_txs_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pcie_ip_txs_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [65:0] pcie_ip_txs_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // pcie_ip_txs_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pcie_ip_txs_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pcie_ip_txs_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // pcie_ip_txs_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pcie_ip_txs_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                      // sdram_s1_translator:uav_waitrequest -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                       // sdram_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_s1_translator:uav_burstcount
	wire   [31:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                        // sdram_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_s1_translator:uav_writedata
	wire   [31:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                          // sdram_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_s1_translator:uav_address
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                            // sdram_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_s1_translator:uav_write
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                             // sdram_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_s1_translator:uav_lock
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                             // sdram_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_s1_translator:uav_read
	wire   [31:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                         // sdram_s1_translator:uav_readdata -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                    // sdram_s1_translator:uav_readdatavalid -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                      // sdram_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_s1_translator:uav_debugaccess
	wire    [3:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                       // sdram_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_s1_translator:uav_byteenable
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                               // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                     // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                             // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                      // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                     // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                            // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                  // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                          // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                   // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                  // sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                 // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                // sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                // sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                 // sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          pcie_ip_bar1_0_translator_avalon_universal_master_0_waitrequest;                                        // pcie_ip_bar1_0_translator_avalon_universal_master_0_agent:av_waitrequest -> pcie_ip_bar1_0_translator:uav_waitrequest
	wire    [9:0] pcie_ip_bar1_0_translator_avalon_universal_master_0_burstcount;                                         // pcie_ip_bar1_0_translator:uav_burstcount -> pcie_ip_bar1_0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [63:0] pcie_ip_bar1_0_translator_avalon_universal_master_0_writedata;                                          // pcie_ip_bar1_0_translator:uav_writedata -> pcie_ip_bar1_0_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] pcie_ip_bar1_0_translator_avalon_universal_master_0_address;                                            // pcie_ip_bar1_0_translator:uav_address -> pcie_ip_bar1_0_translator_avalon_universal_master_0_agent:av_address
	wire          pcie_ip_bar1_0_translator_avalon_universal_master_0_lock;                                               // pcie_ip_bar1_0_translator:uav_lock -> pcie_ip_bar1_0_translator_avalon_universal_master_0_agent:av_lock
	wire          pcie_ip_bar1_0_translator_avalon_universal_master_0_write;                                              // pcie_ip_bar1_0_translator:uav_write -> pcie_ip_bar1_0_translator_avalon_universal_master_0_agent:av_write
	wire          pcie_ip_bar1_0_translator_avalon_universal_master_0_read;                                               // pcie_ip_bar1_0_translator:uav_read -> pcie_ip_bar1_0_translator_avalon_universal_master_0_agent:av_read
	wire   [63:0] pcie_ip_bar1_0_translator_avalon_universal_master_0_readdata;                                           // pcie_ip_bar1_0_translator_avalon_universal_master_0_agent:av_readdata -> pcie_ip_bar1_0_translator:uav_readdata
	wire          pcie_ip_bar1_0_translator_avalon_universal_master_0_debugaccess;                                        // pcie_ip_bar1_0_translator:uav_debugaccess -> pcie_ip_bar1_0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [7:0] pcie_ip_bar1_0_translator_avalon_universal_master_0_byteenable;                                         // pcie_ip_bar1_0_translator:uav_byteenable -> pcie_ip_bar1_0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          pcie_ip_bar1_0_translator_avalon_universal_master_0_readdatavalid;                                      // pcie_ip_bar1_0_translator_avalon_universal_master_0_agent:av_readdatavalid -> pcie_ip_bar1_0_translator:uav_readdatavalid
	wire          custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // custom_slave_block_0_avalon_slave_translator:uav_waitrequest -> custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> custom_slave_block_0_avalon_slave_translator:uav_burstcount
	wire   [31:0] custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> custom_slave_block_0_avalon_slave_translator:uav_writedata
	wire   [31:0] custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_address -> custom_slave_block_0_avalon_slave_translator:uav_address
	wire          custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_write -> custom_slave_block_0_avalon_slave_translator:uav_write
	wire          custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_lock -> custom_slave_block_0_avalon_slave_translator:uav_lock
	wire          custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_read -> custom_slave_block_0_avalon_slave_translator:uav_read
	wire   [31:0] custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // custom_slave_block_0_avalon_slave_translator:uav_readdata -> custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // custom_slave_block_0_avalon_slave_translator:uav_readdatavalid -> custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> custom_slave_block_0_avalon_slave_translator:uav_debugaccess
	wire    [3:0] custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> custom_slave_block_0_avalon_slave_translator:uav_byteenable
	wire          custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [106:0] custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [106:0] custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;       // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;        // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;       // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          pcie_ip_bar2_translator_avalon_universal_master_0_agent_cp_endofpacket;                                 // pcie_ip_bar2_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          pcie_ip_bar2_translator_avalon_universal_master_0_agent_cp_valid;                                       // pcie_ip_bar2_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          pcie_ip_bar2_translator_avalon_universal_master_0_agent_cp_startofpacket;                               // pcie_ip_bar2_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [141:0] pcie_ip_bar2_translator_avalon_universal_master_0_agent_cp_data;                                        // pcie_ip_bar2_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          pcie_ip_bar2_translator_avalon_universal_master_0_agent_cp_ready;                                       // addr_router:sink_ready -> pcie_ip_bar2_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // sgdma_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          sgdma_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                           // sgdma_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          sgdma_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // sgdma_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [105:0] sgdma_csr_translator_avalon_universal_slave_0_agent_rp_data;                                            // sgdma_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          sgdma_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router:sink_ready -> sgdma_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pcie_ip_cra_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // pcie_ip_cra_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          pcie_ip_cra_translator_avalon_universal_slave_0_agent_rp_valid;                                         // pcie_ip_cra_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          pcie_ip_cra_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // pcie_ip_cra_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [105:0] pcie_ip_cra_translator_avalon_universal_slave_0_agent_rp_data;                                          // pcie_ip_cra_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          pcie_ip_cra_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_001:sink_ready -> pcie_ip_cra_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // sgdma_descriptor_read_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid;                              // sgdma_descriptor_read_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // sgdma_descriptor_read_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [108:0] sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_data;                               // sgdma_descriptor_read_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router_001:sink_ready -> sgdma_descriptor_read_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket;                       // sgdma_descriptor_write_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid;                             // sgdma_descriptor_write_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket;                     // sgdma_descriptor_write_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [108:0] sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_data;                              // sgdma_descriptor_write_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready;                             // addr_router_002:sink_ready -> sgdma_descriptor_write_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket;                                 // sgdma_m_read_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire          sgdma_m_read_translator_avalon_universal_master_0_agent_cp_valid;                                       // sgdma_m_read_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire          sgdma_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket;                               // sgdma_m_read_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire  [144:0] sgdma_m_read_translator_avalon_universal_master_0_agent_cp_data;                                        // sgdma_m_read_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire          sgdma_m_read_translator_avalon_universal_master_0_agent_cp_ready;                                       // addr_router_003:sink_ready -> sgdma_m_read_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_m_write_translator_avalon_universal_master_0_agent_cp_endofpacket;                                // sgdma_m_write_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_004:sink_endofpacket
	wire          sgdma_m_write_translator_avalon_universal_master_0_agent_cp_valid;                                      // sgdma_m_write_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_004:sink_valid
	wire          sgdma_m_write_translator_avalon_universal_master_0_agent_cp_startofpacket;                              // sgdma_m_write_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_004:sink_startofpacket
	wire  [144:0] sgdma_m_write_translator_avalon_universal_master_0_agent_cp_data;                                       // sgdma_m_write_translator_avalon_universal_master_0_agent:cp_data -> addr_router_004:sink_data
	wire          sgdma_m_write_translator_avalon_universal_master_0_agent_cp_ready;                                      // addr_router_004:sink_ready -> sgdma_m_write_translator_avalon_universal_master_0_agent:cp_ready
	wire          pcie_ip_txs_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // pcie_ip_txs_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          pcie_ip_txs_translator_avalon_universal_slave_0_agent_rp_valid;                                         // pcie_ip_txs_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          pcie_ip_txs_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // pcie_ip_txs_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [144:0] pcie_ip_txs_translator_avalon_universal_slave_0_agent_rp_data;                                          // pcie_ip_txs_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          pcie_ip_txs_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_002:sink_ready -> pcie_ip_txs_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                      // sdram_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                            // sdram_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                    // sdram_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [108:0] sdram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                             // sdram_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                            // id_router_003:sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pcie_ip_bar1_0_translator_avalon_universal_master_0_agent_cp_endofpacket;                               // pcie_ip_bar1_0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_005:sink_endofpacket
	wire          pcie_ip_bar1_0_translator_avalon_universal_master_0_agent_cp_valid;                                     // pcie_ip_bar1_0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_005:sink_valid
	wire          pcie_ip_bar1_0_translator_avalon_universal_master_0_agent_cp_startofpacket;                             // pcie_ip_bar1_0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_005:sink_startofpacket
	wire  [141:0] pcie_ip_bar1_0_translator_avalon_universal_master_0_agent_cp_data;                                      // pcie_ip_bar1_0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_005:sink_data
	wire          pcie_ip_bar1_0_translator_avalon_universal_master_0_agent_cp_ready;                                     // addr_router_005:sink_ready -> pcie_ip_bar1_0_translator_avalon_universal_master_0_agent:cp_ready
	wire          custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [105:0] custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_004:sink_ready -> custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_src_endofpacket;                                                                            // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                                  // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                                          // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [141:0] addr_router_src_data;                                                                                   // addr_router:src_data -> limiter:cmd_sink_data
	wire    [1:0] addr_router_src_channel;                                                                                // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                                  // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                            // limiter:rsp_src_endofpacket -> pcie_ip_bar2_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                                  // limiter:rsp_src_valid -> pcie_ip_bar2_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                          // limiter:rsp_src_startofpacket -> pcie_ip_bar2_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [141:0] limiter_rsp_src_data;                                                                                   // limiter:rsp_src_data -> pcie_ip_bar2_translator_avalon_universal_master_0_agent:rp_data
	wire    [1:0] limiter_rsp_src_channel;                                                                                // limiter:rsp_src_channel -> pcie_ip_bar2_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                                  // pcie_ip_bar2_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          addr_router_003_src_endofpacket;                                                                        // addr_router_003:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire          addr_router_003_src_valid;                                                                              // addr_router_003:src_valid -> limiter_001:cmd_sink_valid
	wire          addr_router_003_src_startofpacket;                                                                      // addr_router_003:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [144:0] addr_router_003_src_data;                                                                               // addr_router_003:src_data -> limiter_001:cmd_sink_data
	wire    [3:0] addr_router_003_src_channel;                                                                            // addr_router_003:src_channel -> limiter_001:cmd_sink_channel
	wire          addr_router_003_src_ready;                                                                              // limiter_001:cmd_sink_ready -> addr_router_003:src_ready
	wire          limiter_001_rsp_src_endofpacket;                                                                        // limiter_001:rsp_src_endofpacket -> sgdma_m_read_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_001_rsp_src_valid;                                                                              // limiter_001:rsp_src_valid -> sgdma_m_read_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_001_rsp_src_startofpacket;                                                                      // limiter_001:rsp_src_startofpacket -> sgdma_m_read_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [144:0] limiter_001_rsp_src_data;                                                                               // limiter_001:rsp_src_data -> sgdma_m_read_translator_avalon_universal_master_0_agent:rp_data
	wire    [3:0] limiter_001_rsp_src_channel;                                                                            // limiter_001:rsp_src_channel -> sgdma_m_read_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_001_rsp_src_ready;                                                                              // sgdma_m_read_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire          burst_adapter_source0_endofpacket;                                                                      // burst_adapter:source0_endofpacket -> sgdma_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                            // burst_adapter:source0_valid -> sgdma_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                    // burst_adapter:source0_startofpacket -> sgdma_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [105:0] burst_adapter_source0_data;                                                                             // burst_adapter:source0_data -> sgdma_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                            // sgdma_csr_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire    [1:0] burst_adapter_source0_channel;                                                                          // burst_adapter:source0_channel -> sgdma_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_001_source0_endofpacket;                                                                  // burst_adapter_001:source0_endofpacket -> pcie_ip_cra_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_001_source0_valid;                                                                        // burst_adapter_001:source0_valid -> pcie_ip_cra_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_001_source0_startofpacket;                                                                // burst_adapter_001:source0_startofpacket -> pcie_ip_cra_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [105:0] burst_adapter_001_source0_data;                                                                         // burst_adapter_001:source0_data -> pcie_ip_cra_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_001_source0_ready;                                                                        // pcie_ip_cra_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire    [1:0] burst_adapter_001_source0_channel;                                                                      // burst_adapter_001:source0_channel -> pcie_ip_cra_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_002_source0_endofpacket;                                                                  // burst_adapter_002:source0_endofpacket -> pcie_ip_txs_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_002_source0_valid;                                                                        // burst_adapter_002:source0_valid -> pcie_ip_txs_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_002_source0_startofpacket;                                                                // burst_adapter_002:source0_startofpacket -> pcie_ip_txs_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [144:0] burst_adapter_002_source0_data;                                                                         // burst_adapter_002:source0_data -> pcie_ip_txs_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_002_source0_ready;                                                                        // pcie_ip_txs_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_002:source0_ready
	wire    [3:0] burst_adapter_002_source0_channel;                                                                      // burst_adapter_002:source0_channel -> pcie_ip_txs_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_003_source0_endofpacket;                                                                  // burst_adapter_003:source0_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_003_source0_valid;                                                                        // burst_adapter_003:source0_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_003_source0_startofpacket;                                                                // burst_adapter_003:source0_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] burst_adapter_003_source0_data;                                                                         // burst_adapter_003:source0_data -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_003_source0_ready;                                                                        // sdram_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_003:source0_ready
	wire    [3:0] burst_adapter_003_source0_channel;                                                                      // burst_adapter_003:source0_channel -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_004_source0_endofpacket;                                                                  // burst_adapter_004:source0_endofpacket -> custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_004_source0_valid;                                                                        // burst_adapter_004:source0_valid -> custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_004_source0_startofpacket;                                                                // burst_adapter_004:source0_startofpacket -> custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [105:0] burst_adapter_004_source0_data;                                                                         // burst_adapter_004:source0_data -> custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_004_source0_ready;                                                                        // custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_004:source0_ready
	wire    [0:0] burst_adapter_004_source0_channel;                                                                      // burst_adapter_004:source0_channel -> custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                         // rst_controller:reset_out -> [addr_router_001:reset, addr_router_002:reset, addr_router_003:reset, addr_router_004:reset, burst_adapter:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_demux_004:reset, crosser_002:in_reset, crosser_003:in_reset, crosser_004:out_reset, crosser_005:out_reset, id_router:reset, limiter_001:reset, rsp_xbar_demux:reset, rsp_xbar_mux_003:reset, rsp_xbar_mux_004:reset, sgdma:system_reset_n, sgdma_csr_translator:reset, sgdma_csr_translator_avalon_universal_slave_0_agent:reset, sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sgdma_descriptor_read_translator:reset, sgdma_descriptor_read_translator_avalon_universal_master_0_agent:reset, sgdma_descriptor_write_translator:reset, sgdma_descriptor_write_translator_avalon_universal_master_0_agent:reset, sgdma_m_read_translator:reset, sgdma_m_read_translator_avalon_universal_master_0_agent:reset, sgdma_m_write_translator:reset, sgdma_m_write_translator_avalon_universal_master_0_agent:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_004:reset, width_adapter_005:reset, width_adapter_006:reset, width_adapter_007:reset]
	wire          pcie_ip_pcie_core_reset_reset;                                                                          // pcie_ip:pcie_core_reset_reset_n -> [irq_mapper:reset, rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_003:reset_in0]
	wire          rst_controller_001_reset_out_reset;                                                                     // rst_controller_001:reset_out -> [altpll_qsys:reset, burst_adapter_003:reset, cmd_xbar_mux_003:reset, crosser_002:out_reset, crosser_003:out_reset, crosser_004:in_reset, crosser_005:in_reset, id_router_003:reset, rsp_xbar_demux_003:reset, sdram:reset_n, sdram_s1_translator:reset, sdram_s1_translator_avalon_universal_slave_0_agent:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter_010:reset, width_adapter_011:reset]
	wire          rst_controller_002_reset_out_reset;                                                                     // rst_controller_002:reset_out -> [burst_adapter_004:reset, crosser:out_reset, crosser_001:in_reset, custom_slave_block_0:reset_n, custom_slave_block_0_avalon_slave_translator:reset, custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent:reset, custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_004:reset, rsp_xbar_demux_004:reset, width_adapter_012:reset, width_adapter_013:reset]
	wire          rst_controller_003_reset_out_reset;                                                                     // rst_controller_003:reset_out -> [addr_router:reset, addr_router_005:reset, burst_adapter_001:reset, burst_adapter_002:reset, cmd_xbar_demux:reset, cmd_xbar_demux_005:reset, cmd_xbar_mux_002:reset, crosser:in_reset, crosser_001:out_reset, id_router_001:reset, id_router_002:reset, limiter:reset, pcie_ip_bar1_0_translator:reset, pcie_ip_bar1_0_translator_avalon_universal_master_0_agent:reset, pcie_ip_bar2_translator:reset, pcie_ip_bar2_translator_avalon_universal_master_0_agent:reset, pcie_ip_cra_translator:reset, pcie_ip_cra_translator_avalon_universal_slave_0_agent:reset, pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pcie_ip_txs_translator:reset, pcie_ip_txs_translator_avalon_universal_slave_0_agent:reset, pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_mux:reset, width_adapter_002:reset, width_adapter_003:reset, width_adapter_008:reset, width_adapter_009:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                        // cmd_xbar_demux:src0_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                              // cmd_xbar_demux:src0_valid -> width_adapter:in_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                      // cmd_xbar_demux:src0_startofpacket -> width_adapter:in_startofpacket
	wire  [141:0] cmd_xbar_demux_src0_data;                                                                               // cmd_xbar_demux:src0_data -> width_adapter:in_data
	wire    [1:0] cmd_xbar_demux_src0_channel;                                                                            // cmd_xbar_demux:src0_channel -> width_adapter:in_channel
	wire          cmd_xbar_demux_src1_endofpacket;                                                                        // cmd_xbar_demux:src1_endofpacket -> width_adapter_002:in_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                              // cmd_xbar_demux:src1_valid -> width_adapter_002:in_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                      // cmd_xbar_demux:src1_startofpacket -> width_adapter_002:in_startofpacket
	wire  [141:0] cmd_xbar_demux_src1_data;                                                                               // cmd_xbar_demux:src1_data -> width_adapter_002:in_data
	wire    [1:0] cmd_xbar_demux_src1_channel;                                                                            // cmd_xbar_demux:src1_channel -> width_adapter_002:in_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                                                        // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                              // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                      // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [141:0] rsp_xbar_demux_src0_data;                                                                               // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire    [1:0] rsp_xbar_demux_src0_channel;                                                                            // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                              // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                    // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                          // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                                  // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [141:0] rsp_xbar_demux_001_src0_data;                                                                           // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire    [1:0] rsp_xbar_demux_001_src0_channel;                                                                        // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                          // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          limiter_cmd_src_endofpacket;                                                                            // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                                          // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [141:0] limiter_cmd_src_data;                                                                                   // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire    [1:0] limiter_cmd_src_channel;                                                                                // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_cmd_src_ready;                                                                                  // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                           // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                                 // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                         // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [141:0] rsp_xbar_mux_src_data;                                                                                  // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire    [1:0] rsp_xbar_mux_src_channel;                                                                               // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_src_ready;                                                                                 // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire          cmd_xbar_demux_003_src0_endofpacket;                                                                    // cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_002:sink2_endofpacket
	wire          cmd_xbar_demux_003_src0_valid;                                                                          // cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_002:sink2_valid
	wire          cmd_xbar_demux_003_src0_startofpacket;                                                                  // cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_002:sink2_startofpacket
	wire  [144:0] cmd_xbar_demux_003_src0_data;                                                                           // cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_002:sink2_data
	wire    [3:0] cmd_xbar_demux_003_src0_channel;                                                                        // cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_002:sink2_channel
	wire          cmd_xbar_demux_003_src0_ready;                                                                          // cmd_xbar_mux_002:sink2_ready -> cmd_xbar_demux_003:src0_ready
	wire          cmd_xbar_demux_004_src0_endofpacket;                                                                    // cmd_xbar_demux_004:src0_endofpacket -> cmd_xbar_mux_002:sink3_endofpacket
	wire          cmd_xbar_demux_004_src0_valid;                                                                          // cmd_xbar_demux_004:src0_valid -> cmd_xbar_mux_002:sink3_valid
	wire          cmd_xbar_demux_004_src0_startofpacket;                                                                  // cmd_xbar_demux_004:src0_startofpacket -> cmd_xbar_mux_002:sink3_startofpacket
	wire  [144:0] cmd_xbar_demux_004_src0_data;                                                                           // cmd_xbar_demux_004:src0_data -> cmd_xbar_mux_002:sink3_data
	wire    [3:0] cmd_xbar_demux_004_src0_channel;                                                                        // cmd_xbar_demux_004:src0_channel -> cmd_xbar_mux_002:sink3_channel
	wire          cmd_xbar_demux_004_src0_ready;                                                                          // cmd_xbar_mux_002:sink3_ready -> cmd_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_002_src2_endofpacket;                                                                    // rsp_xbar_demux_002:src2_endofpacket -> rsp_xbar_mux_003:sink0_endofpacket
	wire          rsp_xbar_demux_002_src2_valid;                                                                          // rsp_xbar_demux_002:src2_valid -> rsp_xbar_mux_003:sink0_valid
	wire          rsp_xbar_demux_002_src2_startofpacket;                                                                  // rsp_xbar_demux_002:src2_startofpacket -> rsp_xbar_mux_003:sink0_startofpacket
	wire  [144:0] rsp_xbar_demux_002_src2_data;                                                                           // rsp_xbar_demux_002:src2_data -> rsp_xbar_mux_003:sink0_data
	wire    [3:0] rsp_xbar_demux_002_src2_channel;                                                                        // rsp_xbar_demux_002:src2_channel -> rsp_xbar_mux_003:sink0_channel
	wire          rsp_xbar_demux_002_src2_ready;                                                                          // rsp_xbar_mux_003:sink0_ready -> rsp_xbar_demux_002:src2_ready
	wire          rsp_xbar_demux_002_src3_endofpacket;                                                                    // rsp_xbar_demux_002:src3_endofpacket -> rsp_xbar_mux_004:sink0_endofpacket
	wire          rsp_xbar_demux_002_src3_valid;                                                                          // rsp_xbar_demux_002:src3_valid -> rsp_xbar_mux_004:sink0_valid
	wire          rsp_xbar_demux_002_src3_startofpacket;                                                                  // rsp_xbar_demux_002:src3_startofpacket -> rsp_xbar_mux_004:sink0_startofpacket
	wire  [144:0] rsp_xbar_demux_002_src3_data;                                                                           // rsp_xbar_demux_002:src3_data -> rsp_xbar_mux_004:sink0_data
	wire    [3:0] rsp_xbar_demux_002_src3_channel;                                                                        // rsp_xbar_demux_002:src3_channel -> rsp_xbar_mux_004:sink0_channel
	wire          rsp_xbar_demux_002_src3_ready;                                                                          // rsp_xbar_mux_004:sink0_ready -> rsp_xbar_demux_002:src3_ready
	wire          addr_router_001_src_endofpacket;                                                                        // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                              // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                                      // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [108:0] addr_router_001_src_data;                                                                               // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire    [3:0] addr_router_001_src_channel;                                                                            // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                              // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          width_adapter_008_src_ready;                                                                            // sgdma_descriptor_read_translator_avalon_universal_master_0_agent:rp_ready -> width_adapter_008:out_ready
	wire          addr_router_002_src_endofpacket;                                                                        // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          addr_router_002_src_valid;                                                                              // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire          addr_router_002_src_startofpacket;                                                                      // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [108:0] addr_router_002_src_data;                                                                               // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire    [3:0] addr_router_002_src_channel;                                                                            // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire          addr_router_002_src_ready;                                                                              // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire          width_adapter_009_src_ready;                                                                            // sgdma_descriptor_write_translator_avalon_universal_master_0_agent:rp_ready -> width_adapter_009:out_ready
	wire          limiter_001_cmd_src_endofpacket;                                                                        // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire          limiter_001_cmd_src_startofpacket;                                                                      // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire  [144:0] limiter_001_cmd_src_data;                                                                               // limiter_001:cmd_src_data -> cmd_xbar_demux_003:sink_data
	wire    [3:0] limiter_001_cmd_src_channel;                                                                            // limiter_001:cmd_src_channel -> cmd_xbar_demux_003:sink_channel
	wire          limiter_001_cmd_src_ready;                                                                              // cmd_xbar_demux_003:sink_ready -> limiter_001:cmd_src_ready
	wire          rsp_xbar_mux_003_src_endofpacket;                                                                       // rsp_xbar_mux_003:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire          rsp_xbar_mux_003_src_valid;                                                                             // rsp_xbar_mux_003:src_valid -> limiter_001:rsp_sink_valid
	wire          rsp_xbar_mux_003_src_startofpacket;                                                                     // rsp_xbar_mux_003:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [144:0] rsp_xbar_mux_003_src_data;                                                                              // rsp_xbar_mux_003:src_data -> limiter_001:rsp_sink_data
	wire    [3:0] rsp_xbar_mux_003_src_channel;                                                                           // rsp_xbar_mux_003:src_channel -> limiter_001:rsp_sink_channel
	wire          rsp_xbar_mux_003_src_ready;                                                                             // limiter_001:rsp_sink_ready -> rsp_xbar_mux_003:src_ready
	wire          addr_router_004_src_endofpacket;                                                                        // addr_router_004:src_endofpacket -> cmd_xbar_demux_004:sink_endofpacket
	wire          addr_router_004_src_valid;                                                                              // addr_router_004:src_valid -> cmd_xbar_demux_004:sink_valid
	wire          addr_router_004_src_startofpacket;                                                                      // addr_router_004:src_startofpacket -> cmd_xbar_demux_004:sink_startofpacket
	wire  [144:0] addr_router_004_src_data;                                                                               // addr_router_004:src_data -> cmd_xbar_demux_004:sink_data
	wire    [3:0] addr_router_004_src_channel;                                                                            // addr_router_004:src_channel -> cmd_xbar_demux_004:sink_channel
	wire          addr_router_004_src_ready;                                                                              // cmd_xbar_demux_004:sink_ready -> addr_router_004:src_ready
	wire          rsp_xbar_mux_004_src_endofpacket;                                                                       // rsp_xbar_mux_004:src_endofpacket -> sgdma_m_write_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_004_src_valid;                                                                             // rsp_xbar_mux_004:src_valid -> sgdma_m_write_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_004_src_startofpacket;                                                                     // rsp_xbar_mux_004:src_startofpacket -> sgdma_m_write_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [144:0] rsp_xbar_mux_004_src_data;                                                                              // rsp_xbar_mux_004:src_data -> sgdma_m_write_translator_avalon_universal_master_0_agent:rp_data
	wire    [3:0] rsp_xbar_mux_004_src_channel;                                                                           // rsp_xbar_mux_004:src_channel -> sgdma_m_write_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_004_src_ready;                                                                             // sgdma_m_write_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_004:src_ready
	wire          cmd_xbar_mux_002_src_endofpacket;                                                                       // cmd_xbar_mux_002:src_endofpacket -> burst_adapter_002:sink0_endofpacket
	wire          cmd_xbar_mux_002_src_valid;                                                                             // cmd_xbar_mux_002:src_valid -> burst_adapter_002:sink0_valid
	wire          cmd_xbar_mux_002_src_startofpacket;                                                                     // cmd_xbar_mux_002:src_startofpacket -> burst_adapter_002:sink0_startofpacket
	wire  [144:0] cmd_xbar_mux_002_src_data;                                                                              // cmd_xbar_mux_002:src_data -> burst_adapter_002:sink0_data
	wire    [3:0] cmd_xbar_mux_002_src_channel;                                                                           // cmd_xbar_mux_002:src_channel -> burst_adapter_002:sink0_channel
	wire          cmd_xbar_mux_002_src_ready;                                                                             // burst_adapter_002:sink0_ready -> cmd_xbar_mux_002:src_ready
	wire          id_router_002_src_endofpacket;                                                                          // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                                // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                        // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [144:0] id_router_002_src_data;                                                                                 // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire    [3:0] id_router_002_src_channel;                                                                              // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                                // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_mux_003_src_endofpacket;                                                                       // cmd_xbar_mux_003:src_endofpacket -> burst_adapter_003:sink0_endofpacket
	wire          cmd_xbar_mux_003_src_valid;                                                                             // cmd_xbar_mux_003:src_valid -> burst_adapter_003:sink0_valid
	wire          cmd_xbar_mux_003_src_startofpacket;                                                                     // cmd_xbar_mux_003:src_startofpacket -> burst_adapter_003:sink0_startofpacket
	wire  [108:0] cmd_xbar_mux_003_src_data;                                                                              // cmd_xbar_mux_003:src_data -> burst_adapter_003:sink0_data
	wire    [3:0] cmd_xbar_mux_003_src_channel;                                                                           // cmd_xbar_mux_003:src_channel -> burst_adapter_003:sink0_channel
	wire          cmd_xbar_mux_003_src_ready;                                                                             // burst_adapter_003:sink0_ready -> cmd_xbar_mux_003:src_ready
	wire          id_router_003_src_endofpacket;                                                                          // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                                // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                        // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [108:0] id_router_003_src_data;                                                                                 // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire    [3:0] id_router_003_src_channel;                                                                              // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                                // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          addr_router_005_src_endofpacket;                                                                        // addr_router_005:src_endofpacket -> cmd_xbar_demux_005:sink_endofpacket
	wire          addr_router_005_src_valid;                                                                              // addr_router_005:src_valid -> cmd_xbar_demux_005:sink_valid
	wire          addr_router_005_src_startofpacket;                                                                      // addr_router_005:src_startofpacket -> cmd_xbar_demux_005:sink_startofpacket
	wire  [141:0] addr_router_005_src_data;                                                                               // addr_router_005:src_data -> cmd_xbar_demux_005:sink_data
	wire    [0:0] addr_router_005_src_channel;                                                                            // addr_router_005:src_channel -> cmd_xbar_demux_005:sink_channel
	wire          addr_router_005_src_ready;                                                                              // cmd_xbar_demux_005:sink_ready -> addr_router_005:src_ready
	wire          crosser_001_out_ready;                                                                                  // pcie_ip_bar1_0_translator_avalon_universal_master_0_agent:rp_ready -> crosser_001:out_ready
	wire          cmd_xbar_demux_src0_ready;                                                                              // width_adapter:in_ready -> cmd_xbar_demux:src0_ready
	wire          width_adapter_src_endofpacket;                                                                          // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                                // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                        // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire  [105:0] width_adapter_src_data;                                                                                 // width_adapter:out_data -> burst_adapter:sink0_data
	wire          width_adapter_src_ready;                                                                                // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire    [1:0] width_adapter_src_channel;                                                                              // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire          id_router_src_endofpacket;                                                                              // id_router:src_endofpacket -> width_adapter_001:in_endofpacket
	wire          id_router_src_valid;                                                                                    // id_router:src_valid -> width_adapter_001:in_valid
	wire          id_router_src_startofpacket;                                                                            // id_router:src_startofpacket -> width_adapter_001:in_startofpacket
	wire  [105:0] id_router_src_data;                                                                                     // id_router:src_data -> width_adapter_001:in_data
	wire    [1:0] id_router_src_channel;                                                                                  // id_router:src_channel -> width_adapter_001:in_channel
	wire          id_router_src_ready;                                                                                    // width_adapter_001:in_ready -> id_router:src_ready
	wire          width_adapter_001_src_endofpacket;                                                                      // width_adapter_001:out_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          width_adapter_001_src_valid;                                                                            // width_adapter_001:out_valid -> rsp_xbar_demux:sink_valid
	wire          width_adapter_001_src_startofpacket;                                                                    // width_adapter_001:out_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [141:0] width_adapter_001_src_data;                                                                             // width_adapter_001:out_data -> rsp_xbar_demux:sink_data
	wire          width_adapter_001_src_ready;                                                                            // rsp_xbar_demux:sink_ready -> width_adapter_001:out_ready
	wire    [1:0] width_adapter_001_src_channel;                                                                          // width_adapter_001:out_channel -> rsp_xbar_demux:sink_channel
	wire          cmd_xbar_demux_src1_ready;                                                                              // width_adapter_002:in_ready -> cmd_xbar_demux:src1_ready
	wire          width_adapter_002_src_endofpacket;                                                                      // width_adapter_002:out_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire          width_adapter_002_src_valid;                                                                            // width_adapter_002:out_valid -> burst_adapter_001:sink0_valid
	wire          width_adapter_002_src_startofpacket;                                                                    // width_adapter_002:out_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire  [105:0] width_adapter_002_src_data;                                                                             // width_adapter_002:out_data -> burst_adapter_001:sink0_data
	wire          width_adapter_002_src_ready;                                                                            // burst_adapter_001:sink0_ready -> width_adapter_002:out_ready
	wire    [1:0] width_adapter_002_src_channel;                                                                          // width_adapter_002:out_channel -> burst_adapter_001:sink0_channel
	wire          id_router_001_src_endofpacket;                                                                          // id_router_001:src_endofpacket -> width_adapter_003:in_endofpacket
	wire          id_router_001_src_valid;                                                                                // id_router_001:src_valid -> width_adapter_003:in_valid
	wire          id_router_001_src_startofpacket;                                                                        // id_router_001:src_startofpacket -> width_adapter_003:in_startofpacket
	wire  [105:0] id_router_001_src_data;                                                                                 // id_router_001:src_data -> width_adapter_003:in_data
	wire    [1:0] id_router_001_src_channel;                                                                              // id_router_001:src_channel -> width_adapter_003:in_channel
	wire          id_router_001_src_ready;                                                                                // width_adapter_003:in_ready -> id_router_001:src_ready
	wire          width_adapter_003_src_endofpacket;                                                                      // width_adapter_003:out_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          width_adapter_003_src_valid;                                                                            // width_adapter_003:out_valid -> rsp_xbar_demux_001:sink_valid
	wire          width_adapter_003_src_startofpacket;                                                                    // width_adapter_003:out_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [141:0] width_adapter_003_src_data;                                                                             // width_adapter_003:out_data -> rsp_xbar_demux_001:sink_data
	wire          width_adapter_003_src_ready;                                                                            // rsp_xbar_demux_001:sink_ready -> width_adapter_003:out_ready
	wire    [1:0] width_adapter_003_src_channel;                                                                          // width_adapter_003:out_channel -> rsp_xbar_demux_001:sink_channel
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                    // cmd_xbar_demux_001:src0_endofpacket -> width_adapter_004:in_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                          // cmd_xbar_demux_001:src0_valid -> width_adapter_004:in_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                                  // cmd_xbar_demux_001:src0_startofpacket -> width_adapter_004:in_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src0_data;                                                                           // cmd_xbar_demux_001:src0_data -> width_adapter_004:in_data
	wire    [3:0] cmd_xbar_demux_001_src0_channel;                                                                        // cmd_xbar_demux_001:src0_channel -> width_adapter_004:in_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                          // width_adapter_004:in_ready -> cmd_xbar_demux_001:src0_ready
	wire          width_adapter_004_src_endofpacket;                                                                      // width_adapter_004:out_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire          width_adapter_004_src_valid;                                                                            // width_adapter_004:out_valid -> cmd_xbar_mux_002:sink0_valid
	wire          width_adapter_004_src_startofpacket;                                                                    // width_adapter_004:out_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [144:0] width_adapter_004_src_data;                                                                             // width_adapter_004:out_data -> cmd_xbar_mux_002:sink0_data
	wire          width_adapter_004_src_ready;                                                                            // cmd_xbar_mux_002:sink0_ready -> width_adapter_004:out_ready
	wire    [3:0] width_adapter_004_src_channel;                                                                          // width_adapter_004:out_channel -> cmd_xbar_mux_002:sink0_channel
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                                    // cmd_xbar_demux_002:src0_endofpacket -> width_adapter_005:in_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                          // cmd_xbar_demux_002:src0_valid -> width_adapter_005:in_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                                  // cmd_xbar_demux_002:src0_startofpacket -> width_adapter_005:in_startofpacket
	wire  [108:0] cmd_xbar_demux_002_src0_data;                                                                           // cmd_xbar_demux_002:src0_data -> width_adapter_005:in_data
	wire    [3:0] cmd_xbar_demux_002_src0_channel;                                                                        // cmd_xbar_demux_002:src0_channel -> width_adapter_005:in_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                          // width_adapter_005:in_ready -> cmd_xbar_demux_002:src0_ready
	wire          width_adapter_005_src_endofpacket;                                                                      // width_adapter_005:out_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire          width_adapter_005_src_valid;                                                                            // width_adapter_005:out_valid -> cmd_xbar_mux_002:sink1_valid
	wire          width_adapter_005_src_startofpacket;                                                                    // width_adapter_005:out_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [144:0] width_adapter_005_src_data;                                                                             // width_adapter_005:out_data -> cmd_xbar_mux_002:sink1_data
	wire          width_adapter_005_src_ready;                                                                            // cmd_xbar_mux_002:sink1_ready -> width_adapter_005:out_ready
	wire    [3:0] width_adapter_005_src_channel;                                                                          // width_adapter_005:out_channel -> cmd_xbar_mux_002:sink1_channel
	wire          cmd_xbar_demux_003_src1_endofpacket;                                                                    // cmd_xbar_demux_003:src1_endofpacket -> width_adapter_006:in_endofpacket
	wire          cmd_xbar_demux_003_src1_valid;                                                                          // cmd_xbar_demux_003:src1_valid -> width_adapter_006:in_valid
	wire          cmd_xbar_demux_003_src1_startofpacket;                                                                  // cmd_xbar_demux_003:src1_startofpacket -> width_adapter_006:in_startofpacket
	wire  [144:0] cmd_xbar_demux_003_src1_data;                                                                           // cmd_xbar_demux_003:src1_data -> width_adapter_006:in_data
	wire    [3:0] cmd_xbar_demux_003_src1_channel;                                                                        // cmd_xbar_demux_003:src1_channel -> width_adapter_006:in_channel
	wire          cmd_xbar_demux_003_src1_ready;                                                                          // width_adapter_006:in_ready -> cmd_xbar_demux_003:src1_ready
	wire          cmd_xbar_demux_004_src1_endofpacket;                                                                    // cmd_xbar_demux_004:src1_endofpacket -> width_adapter_007:in_endofpacket
	wire          cmd_xbar_demux_004_src1_valid;                                                                          // cmd_xbar_demux_004:src1_valid -> width_adapter_007:in_valid
	wire          cmd_xbar_demux_004_src1_startofpacket;                                                                  // cmd_xbar_demux_004:src1_startofpacket -> width_adapter_007:in_startofpacket
	wire  [144:0] cmd_xbar_demux_004_src1_data;                                                                           // cmd_xbar_demux_004:src1_data -> width_adapter_007:in_data
	wire    [3:0] cmd_xbar_demux_004_src1_channel;                                                                        // cmd_xbar_demux_004:src1_channel -> width_adapter_007:in_channel
	wire          cmd_xbar_demux_004_src1_ready;                                                                          // width_adapter_007:in_ready -> cmd_xbar_demux_004:src1_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                    // rsp_xbar_demux_002:src0_endofpacket -> width_adapter_008:in_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                          // rsp_xbar_demux_002:src0_valid -> width_adapter_008:in_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                                  // rsp_xbar_demux_002:src0_startofpacket -> width_adapter_008:in_startofpacket
	wire  [144:0] rsp_xbar_demux_002_src0_data;                                                                           // rsp_xbar_demux_002:src0_data -> width_adapter_008:in_data
	wire    [3:0] rsp_xbar_demux_002_src0_channel;                                                                        // rsp_xbar_demux_002:src0_channel -> width_adapter_008:in_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                          // width_adapter_008:in_ready -> rsp_xbar_demux_002:src0_ready
	wire          width_adapter_008_src_endofpacket;                                                                      // width_adapter_008:out_endofpacket -> sgdma_descriptor_read_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          width_adapter_008_src_valid;                                                                            // width_adapter_008:out_valid -> sgdma_descriptor_read_translator_avalon_universal_master_0_agent:rp_valid
	wire          width_adapter_008_src_startofpacket;                                                                    // width_adapter_008:out_startofpacket -> sgdma_descriptor_read_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [108:0] width_adapter_008_src_data;                                                                             // width_adapter_008:out_data -> sgdma_descriptor_read_translator_avalon_universal_master_0_agent:rp_data
	wire    [3:0] width_adapter_008_src_channel;                                                                          // width_adapter_008:out_channel -> sgdma_descriptor_read_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_002_src1_endofpacket;                                                                    // rsp_xbar_demux_002:src1_endofpacket -> width_adapter_009:in_endofpacket
	wire          rsp_xbar_demux_002_src1_valid;                                                                          // rsp_xbar_demux_002:src1_valid -> width_adapter_009:in_valid
	wire          rsp_xbar_demux_002_src1_startofpacket;                                                                  // rsp_xbar_demux_002:src1_startofpacket -> width_adapter_009:in_startofpacket
	wire  [144:0] rsp_xbar_demux_002_src1_data;                                                                           // rsp_xbar_demux_002:src1_data -> width_adapter_009:in_data
	wire    [3:0] rsp_xbar_demux_002_src1_channel;                                                                        // rsp_xbar_demux_002:src1_channel -> width_adapter_009:in_channel
	wire          rsp_xbar_demux_002_src1_ready;                                                                          // width_adapter_009:in_ready -> rsp_xbar_demux_002:src1_ready
	wire          width_adapter_009_src_endofpacket;                                                                      // width_adapter_009:out_endofpacket -> sgdma_descriptor_write_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          width_adapter_009_src_valid;                                                                            // width_adapter_009:out_valid -> sgdma_descriptor_write_translator_avalon_universal_master_0_agent:rp_valid
	wire          width_adapter_009_src_startofpacket;                                                                    // width_adapter_009:out_startofpacket -> sgdma_descriptor_write_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [108:0] width_adapter_009_src_data;                                                                             // width_adapter_009:out_data -> sgdma_descriptor_write_translator_avalon_universal_master_0_agent:rp_data
	wire    [3:0] width_adapter_009_src_channel;                                                                          // width_adapter_009:out_channel -> sgdma_descriptor_write_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                    // rsp_xbar_demux_003:src0_endofpacket -> width_adapter_010:in_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                          // rsp_xbar_demux_003:src0_valid -> width_adapter_010:in_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                                  // rsp_xbar_demux_003:src0_startofpacket -> width_adapter_010:in_startofpacket
	wire  [108:0] rsp_xbar_demux_003_src0_data;                                                                           // rsp_xbar_demux_003:src0_data -> width_adapter_010:in_data
	wire    [3:0] rsp_xbar_demux_003_src0_channel;                                                                        // rsp_xbar_demux_003:src0_channel -> width_adapter_010:in_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                          // width_adapter_010:in_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_003_src1_endofpacket;                                                                    // rsp_xbar_demux_003:src1_endofpacket -> width_adapter_011:in_endofpacket
	wire          rsp_xbar_demux_003_src1_valid;                                                                          // rsp_xbar_demux_003:src1_valid -> width_adapter_011:in_valid
	wire          rsp_xbar_demux_003_src1_startofpacket;                                                                  // rsp_xbar_demux_003:src1_startofpacket -> width_adapter_011:in_startofpacket
	wire  [108:0] rsp_xbar_demux_003_src1_data;                                                                           // rsp_xbar_demux_003:src1_data -> width_adapter_011:in_data
	wire    [3:0] rsp_xbar_demux_003_src1_channel;                                                                        // rsp_xbar_demux_003:src1_channel -> width_adapter_011:in_channel
	wire          rsp_xbar_demux_003_src1_ready;                                                                          // width_adapter_011:in_ready -> rsp_xbar_demux_003:src1_ready
	wire          crosser_out_ready;                                                                                      // width_adapter_012:in_ready -> crosser:out_ready
	wire          width_adapter_012_src_endofpacket;                                                                      // width_adapter_012:out_endofpacket -> burst_adapter_004:sink0_endofpacket
	wire          width_adapter_012_src_valid;                                                                            // width_adapter_012:out_valid -> burst_adapter_004:sink0_valid
	wire          width_adapter_012_src_startofpacket;                                                                    // width_adapter_012:out_startofpacket -> burst_adapter_004:sink0_startofpacket
	wire  [105:0] width_adapter_012_src_data;                                                                             // width_adapter_012:out_data -> burst_adapter_004:sink0_data
	wire          width_adapter_012_src_ready;                                                                            // burst_adapter_004:sink0_ready -> width_adapter_012:out_ready
	wire    [0:0] width_adapter_012_src_channel;                                                                          // width_adapter_012:out_channel -> burst_adapter_004:sink0_channel
	wire          id_router_004_src_endofpacket;                                                                          // id_router_004:src_endofpacket -> width_adapter_013:in_endofpacket
	wire          id_router_004_src_valid;                                                                                // id_router_004:src_valid -> width_adapter_013:in_valid
	wire          id_router_004_src_startofpacket;                                                                        // id_router_004:src_startofpacket -> width_adapter_013:in_startofpacket
	wire  [105:0] id_router_004_src_data;                                                                                 // id_router_004:src_data -> width_adapter_013:in_data
	wire    [0:0] id_router_004_src_channel;                                                                              // id_router_004:src_channel -> width_adapter_013:in_channel
	wire          id_router_004_src_ready;                                                                                // width_adapter_013:in_ready -> id_router_004:src_ready
	wire          width_adapter_013_src_endofpacket;                                                                      // width_adapter_013:out_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          width_adapter_013_src_valid;                                                                            // width_adapter_013:out_valid -> rsp_xbar_demux_004:sink_valid
	wire          width_adapter_013_src_startofpacket;                                                                    // width_adapter_013:out_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [141:0] width_adapter_013_src_data;                                                                             // width_adapter_013:out_data -> rsp_xbar_demux_004:sink_data
	wire          width_adapter_013_src_ready;                                                                            // rsp_xbar_demux_004:sink_ready -> width_adapter_013:out_ready
	wire    [0:0] width_adapter_013_src_channel;                                                                          // width_adapter_013:out_channel -> rsp_xbar_demux_004:sink_channel
	wire          crosser_out_endofpacket;                                                                                // crosser:out_endofpacket -> width_adapter_012:in_endofpacket
	wire          crosser_out_valid;                                                                                      // crosser:out_valid -> width_adapter_012:in_valid
	wire          crosser_out_startofpacket;                                                                              // crosser:out_startofpacket -> width_adapter_012:in_startofpacket
	wire  [141:0] crosser_out_data;                                                                                       // crosser:out_data -> width_adapter_012:in_data
	wire          crosser_out_channel;                                                                                    // crosser:out_channel -> width_adapter_012:in_channel
	wire          cmd_xbar_demux_005_src0_endofpacket;                                                                    // cmd_xbar_demux_005:src0_endofpacket -> crosser:in_endofpacket
	wire          cmd_xbar_demux_005_src0_valid;                                                                          // cmd_xbar_demux_005:src0_valid -> crosser:in_valid
	wire          cmd_xbar_demux_005_src0_startofpacket;                                                                  // cmd_xbar_demux_005:src0_startofpacket -> crosser:in_startofpacket
	wire  [141:0] cmd_xbar_demux_005_src0_data;                                                                           // cmd_xbar_demux_005:src0_data -> crosser:in_data
	wire    [0:0] cmd_xbar_demux_005_src0_channel;                                                                        // cmd_xbar_demux_005:src0_channel -> crosser:in_channel
	wire          cmd_xbar_demux_005_src0_ready;                                                                          // crosser:in_ready -> cmd_xbar_demux_005:src0_ready
	wire          crosser_001_out_endofpacket;                                                                            // crosser_001:out_endofpacket -> pcie_ip_bar1_0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          crosser_001_out_valid;                                                                                  // crosser_001:out_valid -> pcie_ip_bar1_0_translator_avalon_universal_master_0_agent:rp_valid
	wire          crosser_001_out_startofpacket;                                                                          // crosser_001:out_startofpacket -> pcie_ip_bar1_0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [141:0] crosser_001_out_data;                                                                                   // crosser_001:out_data -> pcie_ip_bar1_0_translator_avalon_universal_master_0_agent:rp_data
	wire          crosser_001_out_channel;                                                                                // crosser_001:out_channel -> pcie_ip_bar1_0_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                    // rsp_xbar_demux_004:src0_endofpacket -> crosser_001:in_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                          // rsp_xbar_demux_004:src0_valid -> crosser_001:in_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                                  // rsp_xbar_demux_004:src0_startofpacket -> crosser_001:in_startofpacket
	wire  [141:0] rsp_xbar_demux_004_src0_data;                                                                           // rsp_xbar_demux_004:src0_data -> crosser_001:in_data
	wire    [0:0] rsp_xbar_demux_004_src0_channel;                                                                        // rsp_xbar_demux_004:src0_channel -> crosser_001:in_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                          // crosser_001:in_ready -> rsp_xbar_demux_004:src0_ready
	wire          crosser_002_out_endofpacket;                                                                            // crosser_002:out_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire          crosser_002_out_valid;                                                                                  // crosser_002:out_valid -> cmd_xbar_mux_003:sink0_valid
	wire          crosser_002_out_startofpacket;                                                                          // crosser_002:out_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [108:0] crosser_002_out_data;                                                                                   // crosser_002:out_data -> cmd_xbar_mux_003:sink0_data
	wire    [3:0] crosser_002_out_channel;                                                                                // crosser_002:out_channel -> cmd_xbar_mux_003:sink0_channel
	wire          crosser_002_out_ready;                                                                                  // cmd_xbar_mux_003:sink0_ready -> crosser_002:out_ready
	wire          width_adapter_006_src_endofpacket;                                                                      // width_adapter_006:out_endofpacket -> crosser_002:in_endofpacket
	wire          width_adapter_006_src_valid;                                                                            // width_adapter_006:out_valid -> crosser_002:in_valid
	wire          width_adapter_006_src_startofpacket;                                                                    // width_adapter_006:out_startofpacket -> crosser_002:in_startofpacket
	wire  [108:0] width_adapter_006_src_data;                                                                             // width_adapter_006:out_data -> crosser_002:in_data
	wire          width_adapter_006_src_ready;                                                                            // crosser_002:in_ready -> width_adapter_006:out_ready
	wire    [3:0] width_adapter_006_src_channel;                                                                          // width_adapter_006:out_channel -> crosser_002:in_channel
	wire          crosser_003_out_endofpacket;                                                                            // crosser_003:out_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire          crosser_003_out_valid;                                                                                  // crosser_003:out_valid -> cmd_xbar_mux_003:sink1_valid
	wire          crosser_003_out_startofpacket;                                                                          // crosser_003:out_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [108:0] crosser_003_out_data;                                                                                   // crosser_003:out_data -> cmd_xbar_mux_003:sink1_data
	wire    [3:0] crosser_003_out_channel;                                                                                // crosser_003:out_channel -> cmd_xbar_mux_003:sink1_channel
	wire          crosser_003_out_ready;                                                                                  // cmd_xbar_mux_003:sink1_ready -> crosser_003:out_ready
	wire          width_adapter_007_src_endofpacket;                                                                      // width_adapter_007:out_endofpacket -> crosser_003:in_endofpacket
	wire          width_adapter_007_src_valid;                                                                            // width_adapter_007:out_valid -> crosser_003:in_valid
	wire          width_adapter_007_src_startofpacket;                                                                    // width_adapter_007:out_startofpacket -> crosser_003:in_startofpacket
	wire  [108:0] width_adapter_007_src_data;                                                                             // width_adapter_007:out_data -> crosser_003:in_data
	wire          width_adapter_007_src_ready;                                                                            // crosser_003:in_ready -> width_adapter_007:out_ready
	wire    [3:0] width_adapter_007_src_channel;                                                                          // width_adapter_007:out_channel -> crosser_003:in_channel
	wire          crosser_004_out_endofpacket;                                                                            // crosser_004:out_endofpacket -> rsp_xbar_mux_003:sink1_endofpacket
	wire          crosser_004_out_valid;                                                                                  // crosser_004:out_valid -> rsp_xbar_mux_003:sink1_valid
	wire          crosser_004_out_startofpacket;                                                                          // crosser_004:out_startofpacket -> rsp_xbar_mux_003:sink1_startofpacket
	wire  [144:0] crosser_004_out_data;                                                                                   // crosser_004:out_data -> rsp_xbar_mux_003:sink1_data
	wire    [3:0] crosser_004_out_channel;                                                                                // crosser_004:out_channel -> rsp_xbar_mux_003:sink1_channel
	wire          crosser_004_out_ready;                                                                                  // rsp_xbar_mux_003:sink1_ready -> crosser_004:out_ready
	wire          width_adapter_010_src_endofpacket;                                                                      // width_adapter_010:out_endofpacket -> crosser_004:in_endofpacket
	wire          width_adapter_010_src_valid;                                                                            // width_adapter_010:out_valid -> crosser_004:in_valid
	wire          width_adapter_010_src_startofpacket;                                                                    // width_adapter_010:out_startofpacket -> crosser_004:in_startofpacket
	wire  [144:0] width_adapter_010_src_data;                                                                             // width_adapter_010:out_data -> crosser_004:in_data
	wire          width_adapter_010_src_ready;                                                                            // crosser_004:in_ready -> width_adapter_010:out_ready
	wire    [3:0] width_adapter_010_src_channel;                                                                          // width_adapter_010:out_channel -> crosser_004:in_channel
	wire          crosser_005_out_endofpacket;                                                                            // crosser_005:out_endofpacket -> rsp_xbar_mux_004:sink1_endofpacket
	wire          crosser_005_out_valid;                                                                                  // crosser_005:out_valid -> rsp_xbar_mux_004:sink1_valid
	wire          crosser_005_out_startofpacket;                                                                          // crosser_005:out_startofpacket -> rsp_xbar_mux_004:sink1_startofpacket
	wire  [144:0] crosser_005_out_data;                                                                                   // crosser_005:out_data -> rsp_xbar_mux_004:sink1_data
	wire    [3:0] crosser_005_out_channel;                                                                                // crosser_005:out_channel -> rsp_xbar_mux_004:sink1_channel
	wire          crosser_005_out_ready;                                                                                  // rsp_xbar_mux_004:sink1_ready -> crosser_005:out_ready
	wire          width_adapter_011_src_endofpacket;                                                                      // width_adapter_011:out_endofpacket -> crosser_005:in_endofpacket
	wire          width_adapter_011_src_valid;                                                                            // width_adapter_011:out_valid -> crosser_005:in_valid
	wire          width_adapter_011_src_startofpacket;                                                                    // width_adapter_011:out_startofpacket -> crosser_005:in_startofpacket
	wire  [144:0] width_adapter_011_src_data;                                                                             // width_adapter_011:out_data -> crosser_005:in_data
	wire          width_adapter_011_src_ready;                                                                            // crosser_005:in_ready -> width_adapter_011:out_ready
	wire    [3:0] width_adapter_011_src_channel;                                                                          // width_adapter_011:out_channel -> crosser_005:in_channel
	wire    [1:0] limiter_cmd_valid_data;                                                                                 // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire    [3:0] limiter_001_cmd_valid_data;                                                                             // limiter_001:cmd_src_valid -> cmd_xbar_demux_003:sink_valid
	wire          irq_mapper_receiver0_irq;                                                                               // sgdma:csr_irq -> irq_mapper:receiver0_irq
	wire   [15:0] pcie_ip_rxm_irq_irq;                                                                                    // irq_mapper:sender_irq -> pcie_ip:rxm_irq_irq

	amm_master_qsys_with_pcie_pcie_ip #(
		.p_pcie_hip_type                     ("2"),
		.lane_mask                           (8'b11111110),
		.max_link_width                      (1),
		.millisecond_cycle_count             ("125000"),
		.enable_gen2_core                    ("false"),
		.gen2_lane_rate_mode                 ("false"),
		.no_soft_reset                       ("false"),
		.core_clk_divider                    (2),
		.enable_ch0_pclk_out                 ("true"),
		.core_clk_source                     ("pclk"),
		.CB_P2A_AVALON_ADDR_B0               (0),
		.bar0_size_mask                      (7),
		.bar0_io_space                       ("false"),
		.bar0_64bit_mem_space                ("true"),
		.bar0_prefetchable                   ("true"),
		.CB_P2A_AVALON_ADDR_B1               (0),
		.bar1_size_mask                      (0),
		.bar1_io_space                       ("false"),
		.bar1_64bit_mem_space                ("true"),
		.bar1_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B2               (0),
		.bar2_size_mask                      (15),
		.bar2_io_space                       ("false"),
		.bar2_64bit_mem_space                ("false"),
		.bar2_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B3               (0),
		.bar3_size_mask                      (0),
		.bar3_io_space                       ("false"),
		.bar3_64bit_mem_space                ("false"),
		.bar3_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B4               (0),
		.bar4_size_mask                      (0),
		.bar4_io_space                       ("false"),
		.bar4_64bit_mem_space                ("false"),
		.bar4_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B5               (0),
		.bar5_size_mask                      (0),
		.bar5_io_space                       ("false"),
		.bar5_64bit_mem_space                ("false"),
		.bar5_prefetchable                   ("false"),
		.vendor_id                           (4466),
		.device_id                           (57345),
		.revision_id                         (1),
		.class_code                          (0),
		.subsystem_vendor_id                 (4466),
		.subsystem_device_id                 (4),
		.port_link_number                    (1),
		.msi_function_count                  (0),
		.enable_msi_64bit_addressing         ("true"),
		.enable_function_msix_support        ("false"),
		.eie_before_nfts_count               (4),
		.enable_completion_timeout_disable   ("false"),
		.completion_timeout                  ("NONE"),
		.enable_adapter_half_rate_mode       ("false"),
		.msix_pba_bir                        (0),
		.msix_pba_offset                     (0),
		.msix_table_bir                      (0),
		.msix_table_offset                   (0),
		.msix_table_size                     (0),
		.use_crc_forwarding                  ("false"),
		.surprise_down_error_support         ("false"),
		.dll_active_report_support           ("false"),
		.bar_io_window_size                  ("32BIT"),
		.bar_prefetchable                    (32),
		.hot_plug_support                    (7'b0000000),
		.no_command_completed                ("true"),
		.slot_power_limit                    (0),
		.slot_power_scale                    (0),
		.slot_number                         (0),
		.enable_slot_register                ("false"),
		.advanced_errors                     ("false"),
		.enable_ecrc_check                   ("false"),
		.enable_ecrc_gen                     ("false"),
		.max_payload_size                    (0),
		.retry_buffer_last_active_address    (255),
		.credit_buffer_allocation_aux        ("ABSOLUTE"),
		.vc0_rx_flow_ctrl_posted_header      (28),
		.vc0_rx_flow_ctrl_posted_data        (198),
		.vc0_rx_flow_ctrl_nonposted_header   (30),
		.vc0_rx_flow_ctrl_nonposted_data     (0),
		.vc0_rx_flow_ctrl_compl_header       (48),
		.vc0_rx_flow_ctrl_compl_data         (256),
		.RX_BUF                              (9),
		.RH_NUM                              (7),
		.G_TAG_NUM0                          (32),
		.endpoint_l0_latency                 (0),
		.endpoint_l1_latency                 (0),
		.enable_l1_aspm                      ("false"),
		.l01_entry_latency                   (31),
		.diffclock_nfts_count                (255),
		.sameclock_nfts_count                (255),
		.l1_exit_latency_sameclock           (7),
		.l1_exit_latency_diffclock           (7),
		.l0_exit_latency_sameclock           (7),
		.l0_exit_latency_diffclock           (7),
		.gen2_diffclock_nfts_count           (255),
		.gen2_sameclock_nfts_count           (255),
		.CG_COMMON_CLOCK_MODE                (1),
		.CB_PCIE_MODE                        (0),
		.AST_LITE                            (0),
		.CB_PCIE_RX_LITE                     (0),
		.CG_RXM_IRQ_NUM                      (16),
		.CG_AVALON_S_ADDR_WIDTH              (20),
		.bypass_tl                           ("false"),
		.CG_IMPL_CRA_AV_SLAVE_PORT           (1),
		.CG_NO_CPL_REORDERING                (0),
		.CG_ENABLE_A2P_INTERRUPT             (0),
		.CG_IRQ_BIT_ENA                      (65535),
		.CB_A2P_ADDR_MAP_IS_FIXED            (1),
		.CB_A2P_ADDR_MAP_NUM_ENTRIES         (1),
		.CB_A2P_ADDR_MAP_PASS_THRU_BITS      (31),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_0_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_0_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_1_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_1_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_2_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_2_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_3_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_3_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_4_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_4_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_5_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_5_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_6_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_6_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_7_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_7_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_8_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_8_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_9_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_9_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_10_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_10_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_11_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_11_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_12_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_12_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_13_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_13_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_14_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_14_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_15_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_15_LOW  (32'b00000000000000000000000000000000),
		.RXM_DATA_WIDTH                      (64),
		.RXM_BEN_WIDTH                       (8),
		.TL_SELECTION                        (1),
		.pcie_mode                           ("SHARED_MODE"),
		.single_rx_detect                    (1),
		.enable_coreclk_out_half_rate        ("false"),
		.low_priority_vc                     (0),
		.link_width                          (1),
		.cyclone4                            (1)
	) pcie_ip (
		.pcie_core_clk_clk                  (pcie_ip_pcie_core_clk_clk),                                //      pcie_core_clk.clk
		.pcie_core_reset_reset_n            (pcie_ip_pcie_core_reset_reset),                            //    pcie_core_reset.reset_n
		.cal_blk_clk_clk                    (altpll_qsys_c3_clk),                                       //        cal_blk_clk.clk
		.txs_address                        (pcie_ip_txs_translator_avalon_anti_slave_0_address),       //                txs.address
		.txs_chipselect                     (pcie_ip_txs_translator_avalon_anti_slave_0_chipselect),    //                   .chipselect
		.txs_byteenable                     (pcie_ip_txs_translator_avalon_anti_slave_0_byteenable),    //                   .byteenable
		.txs_readdata                       (pcie_ip_txs_translator_avalon_anti_slave_0_readdata),      //                   .readdata
		.txs_writedata                      (pcie_ip_txs_translator_avalon_anti_slave_0_writedata),     //                   .writedata
		.txs_read                           (pcie_ip_txs_translator_avalon_anti_slave_0_read),          //                   .read
		.txs_write                          (pcie_ip_txs_translator_avalon_anti_slave_0_write),         //                   .write
		.txs_burstcount                     (pcie_ip_txs_translator_avalon_anti_slave_0_burstcount),    //                   .burstcount
		.txs_readdatavalid                  (pcie_ip_txs_translator_avalon_anti_slave_0_readdatavalid), //                   .readdatavalid
		.txs_waitrequest                    (pcie_ip_txs_translator_avalon_anti_slave_0_waitrequest),   //                   .waitrequest
		.refclk_export                      (pcie_ip_refclk_export),                                    //             refclk.export
		.test_in_test_in                    (pcie_ip_test_in_test_in),                                  //            test_in.test_in
		.pcie_rstn_export                   (pcie_ip_pcie_rstn_export),                                 //          pcie_rstn.export
		.clocks_sim_clk250_export           (pcie_ip_clocks_sim_clk250_export),                         //         clocks_sim.clk250_export
		.clocks_sim_clk500_export           (pcie_ip_clocks_sim_clk500_export),                         //                   .clk500_export
		.clocks_sim_clk125_export           (pcie_ip_clocks_sim_clk125_export),                         //                   .clk125_export
		.reconfig_busy_busy_altgxb_reconfig (pcie_ip_reconfig_busy_busy_altgxb_reconfig),               //      reconfig_busy.busy_altgxb_reconfig
		.pipe_ext_pipe_mode                 (pcie_ip_pipe_ext_pipe_mode),                               //           pipe_ext.pipe_mode
		.pipe_ext_phystatus_ext             (pcie_ip_pipe_ext_phystatus_ext),                           //                   .phystatus_ext
		.pipe_ext_rate_ext                  (pcie_ip_pipe_ext_rate_ext),                                //                   .rate_ext
		.pipe_ext_powerdown_ext             (pcie_ip_pipe_ext_powerdown_ext),                           //                   .powerdown_ext
		.pipe_ext_txdetectrx_ext            (pcie_ip_pipe_ext_txdetectrx_ext),                          //                   .txdetectrx_ext
		.pipe_ext_rxelecidle0_ext           (pcie_ip_pipe_ext_rxelecidle0_ext),                         //                   .rxelecidle0_ext
		.pipe_ext_rxdata0_ext               (pcie_ip_pipe_ext_rxdata0_ext),                             //                   .rxdata0_ext
		.pipe_ext_rxstatus0_ext             (pcie_ip_pipe_ext_rxstatus0_ext),                           //                   .rxstatus0_ext
		.pipe_ext_rxvalid0_ext              (pcie_ip_pipe_ext_rxvalid0_ext),                            //                   .rxvalid0_ext
		.pipe_ext_rxdatak0_ext              (pcie_ip_pipe_ext_rxdatak0_ext),                            //                   .rxdatak0_ext
		.pipe_ext_txdata0_ext               (pcie_ip_pipe_ext_txdata0_ext),                             //                   .txdata0_ext
		.pipe_ext_txdatak0_ext              (pcie_ip_pipe_ext_txdatak0_ext),                            //                   .txdatak0_ext
		.pipe_ext_rxpolarity0_ext           (pcie_ip_pipe_ext_rxpolarity0_ext),                         //                   .rxpolarity0_ext
		.pipe_ext_txcompl0_ext              (pcie_ip_pipe_ext_txcompl0_ext),                            //                   .txcompl0_ext
		.pipe_ext_txelecidle0_ext           (pcie_ip_pipe_ext_txelecidle0_ext),                         //                   .txelecidle0_ext
		.powerdown_pll_powerdown            (pcie_ip_powerdown_pll_powerdown),                          //          powerdown.pll_powerdown
		.powerdown_gxb_powerdown            (pcie_ip_powerdown_gxb_powerdown),                          //                   .gxb_powerdown
		.bar1_0_address                     (pcie_ip_bar1_0_address),                                   //             bar1_0.address
		.bar1_0_read                        (pcie_ip_bar1_0_read),                                      //                   .read
		.bar1_0_waitrequest                 (pcie_ip_bar1_0_waitrequest),                               //                   .waitrequest
		.bar1_0_write                       (pcie_ip_bar1_0_write),                                     //                   .write
		.bar1_0_readdatavalid               (pcie_ip_bar1_0_readdatavalid),                             //                   .readdatavalid
		.bar1_0_readdata                    (pcie_ip_bar1_0_readdata),                                  //                   .readdata
		.bar1_0_writedata                   (pcie_ip_bar1_0_writedata),                                 //                   .writedata
		.bar1_0_burstcount                  (pcie_ip_bar1_0_burstcount),                                //                   .burstcount
		.bar1_0_byteenable                  (pcie_ip_bar1_0_byteenable),                                //                   .byteenable
		.bar2_address                       (pcie_ip_bar2_address),                                     //               bar2.address
		.bar2_read                          (pcie_ip_bar2_read),                                        //                   .read
		.bar2_waitrequest                   (pcie_ip_bar2_waitrequest),                                 //                   .waitrequest
		.bar2_write                         (pcie_ip_bar2_write),                                       //                   .write
		.bar2_readdatavalid                 (pcie_ip_bar2_readdatavalid),                               //                   .readdatavalid
		.bar2_readdata                      (pcie_ip_bar2_readdata),                                    //                   .readdata
		.bar2_writedata                     (pcie_ip_bar2_writedata),                                   //                   .writedata
		.bar2_burstcount                    (pcie_ip_bar2_burstcount),                                  //                   .burstcount
		.bar2_byteenable                    (pcie_ip_bar2_byteenable),                                  //                   .byteenable
		.cra_chipselect                     (pcie_ip_cra_translator_avalon_anti_slave_0_chipselect),    //                cra.chipselect
		.cra_address                        (pcie_ip_cra_translator_avalon_anti_slave_0_address),       //                   .address
		.cra_byteenable                     (pcie_ip_cra_translator_avalon_anti_slave_0_byteenable),    //                   .byteenable
		.cra_read                           (pcie_ip_cra_translator_avalon_anti_slave_0_read),          //                   .read
		.cra_readdata                       (pcie_ip_cra_translator_avalon_anti_slave_0_readdata),      //                   .readdata
		.cra_write                          (pcie_ip_cra_translator_avalon_anti_slave_0_write),         //                   .write
		.cra_writedata                      (pcie_ip_cra_translator_avalon_anti_slave_0_writedata),     //                   .writedata
		.cra_waitrequest                    (pcie_ip_cra_translator_avalon_anti_slave_0_waitrequest),   //                   .waitrequest
		.cra_irq_irq                        (),                                                         //            cra_irq.irq
		.rxm_irq_irq                        (pcie_ip_rxm_irq_irq),                                      //            rxm_irq.irq
		.rx_in_rx_datain_0                  (pcie_ip_rx_in_rx_datain_0),                                //              rx_in.rx_datain_0
		.tx_out_tx_dataout_0                (pcie_ip_tx_out_tx_dataout_0),                              //             tx_out.tx_dataout_0
		.reconfig_togxb_data                (pcie_ip_reconfig_togxb_data),                              //     reconfig_togxb.data
		.reconfig_gxbclk_clk                (altpll_qsys_c3_clk),                                       //    reconfig_gxbclk.clk
		.reconfig_fromgxb_0_data            (pcie_ip_reconfig_fromgxb_0_data),                          // reconfig_fromgxb_0.data
		.fixedclk_clk                       (pcie_ip_pcie_core_clk_clk)                                 //           fixedclk.clk
	);

	amm_master_qsys_with_pcie_sgdma sgdma (
		.clk                           (pcie_ip_pcie_core_clk_clk),                           //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),                     //            reset.reset_n
		.csr_chipselect                (sgdma_csr_translator_avalon_anti_slave_0_chipselect), //              csr.chipselect
		.csr_address                   (sgdma_csr_translator_avalon_anti_slave_0_address),    //                 .address
		.csr_read                      (sgdma_csr_translator_avalon_anti_slave_0_read),       //                 .read
		.csr_write                     (sgdma_csr_translator_avalon_anti_slave_0_write),      //                 .write
		.csr_writedata                 (sgdma_csr_translator_avalon_anti_slave_0_writedata),  //                 .writedata
		.csr_readdata                  (sgdma_csr_translator_avalon_anti_slave_0_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_descriptor_read_readdata),                      //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_descriptor_read_readdatavalid),                 //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_descriptor_read_waitrequest),                   //                 .waitrequest
		.descriptor_read_address       (sgdma_descriptor_read_address),                       //                 .address
		.descriptor_read_read          (sgdma_descriptor_read_read),                          //                 .read
		.descriptor_write_waitrequest  (sgdma_descriptor_write_waitrequest),                  // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_descriptor_write_address),                      //                 .address
		.descriptor_write_write        (sgdma_descriptor_write_write),                        //                 .write
		.descriptor_write_writedata    (sgdma_descriptor_write_writedata),                    //                 .writedata
		.csr_irq                       (irq_mapper_receiver0_irq),                            //          csr_irq.irq
		.m_read_readdata               (sgdma_m_read_readdata),                               //           m_read.readdata
		.m_read_readdatavalid          (sgdma_m_read_readdatavalid),                          //                 .readdatavalid
		.m_read_waitrequest            (sgdma_m_read_waitrequest),                            //                 .waitrequest
		.m_read_address                (sgdma_m_read_address),                                //                 .address
		.m_read_read                   (sgdma_m_read_read),                                   //                 .read
		.m_read_burstcount             (sgdma_m_read_burstcount),                             //                 .burstcount
		.m_write_waitrequest           (sgdma_m_write_waitrequest),                           //          m_write.waitrequest
		.m_write_address               (sgdma_m_write_address),                               //                 .address
		.m_write_write                 (sgdma_m_write_write),                                 //                 .write
		.m_write_writedata             (sgdma_m_write_writedata),                             //                 .writedata
		.m_write_byteenable            (sgdma_m_write_byteenable),                            //                 .byteenable
		.m_write_burstcount            (sgdma_m_write_burstcount)                             //                 .burstcount
	);

	amm_master_qsys_with_pcie_sdram sdram (
		.clk            (clk_clk),                                               //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                   // reset.reset_n
		.az_addr        (sdram_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                                            //  wire.export
		.zs_ba          (sdram_ba),                                              //      .export
		.zs_cas_n       (sdram_cas_n),                                           //      .export
		.zs_cke         (sdram_cke),                                             //      .export
		.zs_cs_n        (sdram_cs_n),                                            //      .export
		.zs_dq          (sdram_dq),                                              //      .export
		.zs_dqm         (sdram_dqm),                                             //      .export
		.zs_ras_n       (sdram_ras_n),                                           //      .export
		.zs_we_n        (sdram_we_n)                                             //      .export
	);

	amm_master_qsys_with_pcie_altpll_qsys altpll_qsys (
		.clk       (clk_clk),                            //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset), // inclk_interface_reset.reset
		.read      (),                                   //             pll_slave.read
		.write     (),                                   //                      .write
		.address   (),                                   //                      .address
		.readdata  (),                                   //                      .readdata
		.writedata (),                                   //                      .writedata
		.c0        (),                                   //                    c0.clk
		.c1        (altpll_sdram_clk),                   //                    c1.clk
		.c2        (),                                   //                    c2.clk
		.c3        (altpll_qsys_c3_clk),                 //                    c3.clk
		.areset    (),                                   //        areset_conduit.export
		.locked    (),                                   //        locked_conduit.export
		.phasedone ()                                    //     phasedone_conduit.export
	);

	custom_slave #(
		.MASTER_ADDRESSWIDTH (28),
		.SLAVE_ADDRESSWIDTH  (5),
		.DATAWIDTH           (32),
		.NUMREGS             (32),
		.REGWIDTH            (32)
	) custom_slave_block_0 (
		.clk                  (clk_clk),                                                                     //         clock.clk
		.reset_n              (~rst_controller_002_reset_out_reset),                                         //         reset.reset_n
		.master_address       (),                                                                            // avalon_master.address
		.master_writedata     (),                                                                            //              .writedata
		.master_write         (),                                                                            //              .write
		.master_read          (),                                                                            //              .read
		.master_readdata      (),                                                                            //              .readdata
		.master_readdatavalid (),                                                                            //              .readdatavalid
		.master_waitrequest   (),                                                                            //              .waitrequest
		.slave_readdata       (custom_slave_block_0_avalon_slave_translator_avalon_anti_slave_0_readdata),   //  avalon_slave.readdata
		.slave_chipselect     (custom_slave_block_0_avalon_slave_translator_avalon_anti_slave_0_chipselect), //              .chipselect
		.slave_read           (custom_slave_block_0_avalon_slave_translator_avalon_anti_slave_0_read),       //              .read
		.slave_write          (custom_slave_block_0_avalon_slave_translator_avalon_anti_slave_0_write),      //              .write
		.slave_writedata      (custom_slave_block_0_avalon_slave_translator_avalon_anti_slave_0_writedata),  //              .writedata
		.slave_address        (custom_slave_block_0_avalon_slave_translator_avalon_anti_slave_0_address),    //              .address
		.rdwr_cntl            (custom_module_conduit_rdwr_cntl),                                             //   conduit_end.export
		.n_action             (custom_module_conduit_n_action),                                              //              .export
		.add_data_sel         (custom_module_conduit_add_data_sel),                                          //              .export
		.rdwr_address         (custom_module_conduit_rdwr_address)                                           //              .export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (64),
		.AV_BURSTCOUNT_W             (7),
		.AV_BYTEENABLE_W             (8),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (10),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (8),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (1),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) pcie_ip_bar2_translator (
		.clk                      (pcie_ip_pcie_core_clk_clk),                                       //                       clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                              //                     reset.reset
		.uav_address              (pcie_ip_bar2_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (pcie_ip_bar2_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (pcie_ip_bar2_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (pcie_ip_bar2_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (pcie_ip_bar2_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (pcie_ip_bar2_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (pcie_ip_bar2_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (pcie_ip_bar2_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (pcie_ip_bar2_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (pcie_ip_bar2_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (pcie_ip_bar2_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (pcie_ip_bar2_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (pcie_ip_bar2_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (pcie_ip_bar2_burstcount),                                         //                          .burstcount
		.av_byteenable            (pcie_ip_bar2_byteenable),                                         //                          .byteenable
		.av_read                  (pcie_ip_bar2_read),                                               //                          .read
		.av_readdata              (pcie_ip_bar2_readdata),                                           //                          .readdata
		.av_readdatavalid         (pcie_ip_bar2_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (pcie_ip_bar2_write),                                              //                          .write
		.av_writedata             (pcie_ip_bar2_writedata),                                          //                          .writedata
		.av_beginbursttransfer    (1'b0),                                                            //               (terminated)
		.av_begintransfer         (1'b0),                                                            //               (terminated)
		.av_chipselect            (1'b0),                                                            //               (terminated)
		.av_lock                  (1'b0),                                                            //               (terminated)
		.av_debugaccess           (1'b0),                                                            //               (terminated)
		.uav_clken                (),                                                                //               (terminated)
		.av_clken                 (1'b1),                                                            //               (terminated)
		.uav_response             (2'b00),                                                           //               (terminated)
		.av_response              (),                                                                //               (terminated)
		.uav_writeresponserequest (),                                                                //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                            //               (terminated)
		.av_writeresponserequest  (1'b0),                                                            //               (terminated)
		.av_writeresponsevalid    ()                                                                 //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (4),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sgdma_csr_translator (
		.clk                      (pcie_ip_pcie_core_clk_clk),                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address              (sgdma_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sgdma_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sgdma_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sgdma_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sgdma_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sgdma_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sgdma_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sgdma_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sgdma_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sgdma_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sgdma_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sgdma_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sgdma_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (sgdma_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (sgdma_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sgdma_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (sgdma_csr_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                     //              (terminated)
		.av_burstcount            (),                                                                     //              (terminated)
		.av_byteenable            (),                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                 //              (terminated)
		.av_waitrequest           (1'b0),                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                     //              (terminated)
		.av_lock                  (),                                                                     //              (terminated)
		.av_clken                 (),                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                 //              (terminated)
		.av_debugaccess           (),                                                                     //              (terminated)
		.av_outputenable          (),                                                                     //              (terminated)
		.uav_response             (),                                                                     //              (terminated)
		.av_response              (2'b00),                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (12),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pcie_ip_cra_translator (
		.clk                      (pcie_ip_pcie_core_clk_clk),                                              //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                     //                    reset.reset
		.uav_address              (pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pcie_ip_cra_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (pcie_ip_cra_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (pcie_ip_cra_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (pcie_ip_cra_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (pcie_ip_cra_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (pcie_ip_cra_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (pcie_ip_cra_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (pcie_ip_cra_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_descriptor_read_translator (
		.clk                      (pcie_ip_pcie_core_clk_clk),                                                //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                           //                     reset.reset
		.uav_address              (sgdma_descriptor_read_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (sgdma_descriptor_read_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (sgdma_descriptor_read_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (sgdma_descriptor_read_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (sgdma_descriptor_read_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (sgdma_descriptor_read_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (sgdma_descriptor_read_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (sgdma_descriptor_read_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (sgdma_descriptor_read_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (sgdma_descriptor_read_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (sgdma_descriptor_read_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (sgdma_descriptor_read_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (sgdma_descriptor_read_waitrequest),                                        //                          .waitrequest
		.av_read                  (sgdma_descriptor_read_read),                                               //                          .read
		.av_readdata              (sgdma_descriptor_read_readdata),                                           //                          .readdata
		.av_readdatavalid         (sgdma_descriptor_read_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount            (1'b1),                                                                     //               (terminated)
		.av_byteenable            (4'b1111),                                                                  //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                     //               (terminated)
		.av_begintransfer         (1'b0),                                                                     //               (terminated)
		.av_chipselect            (1'b0),                                                                     //               (terminated)
		.av_write                 (1'b0),                                                                     //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                     //               (terminated)
		.av_lock                  (1'b0),                                                                     //               (terminated)
		.av_debugaccess           (1'b0),                                                                     //               (terminated)
		.uav_clken                (),                                                                         //               (terminated)
		.av_clken                 (1'b1),                                                                     //               (terminated)
		.uav_response             (2'b00),                                                                    //               (terminated)
		.av_response              (),                                                                         //               (terminated)
		.uav_writeresponserequest (),                                                                         //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                     //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                     //               (terminated)
		.av_writeresponsevalid    ()                                                                          //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_descriptor_write_translator (
		.clk                      (pcie_ip_pcie_core_clk_clk),                                                 //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                            //                     reset.reset
		.uav_address              (sgdma_descriptor_write_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (sgdma_descriptor_write_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (sgdma_descriptor_write_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (sgdma_descriptor_write_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (sgdma_descriptor_write_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (sgdma_descriptor_write_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (sgdma_descriptor_write_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (sgdma_descriptor_write_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (sgdma_descriptor_write_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (sgdma_descriptor_write_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (sgdma_descriptor_write_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (sgdma_descriptor_write_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (sgdma_descriptor_write_waitrequest),                                        //                          .waitrequest
		.av_write                 (sgdma_descriptor_write_write),                                              //                          .write
		.av_writedata             (sgdma_descriptor_write_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                      //               (terminated)
		.av_byteenable            (4'b1111),                                                                   //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                      //               (terminated)
		.av_begintransfer         (1'b0),                                                                      //               (terminated)
		.av_chipselect            (1'b0),                                                                      //               (terminated)
		.av_read                  (1'b0),                                                                      //               (terminated)
		.av_readdata              (),                                                                          //               (terminated)
		.av_readdatavalid         (),                                                                          //               (terminated)
		.av_lock                  (1'b0),                                                                      //               (terminated)
		.av_debugaccess           (1'b0),                                                                      //               (terminated)
		.uav_clken                (),                                                                          //               (terminated)
		.av_clken                 (1'b1),                                                                      //               (terminated)
		.uav_response             (2'b00),                                                                     //               (terminated)
		.av_response              (),                                                                          //               (terminated)
		.uav_writeresponserequest (),                                                                          //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                      //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                      //               (terminated)
		.av_writeresponsevalid    ()                                                                           //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (64),
		.AV_BURSTCOUNT_W             (4),
		.AV_BYTEENABLE_W             (8),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (7),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (8),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (1),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_m_read_translator (
		.clk                      (pcie_ip_pcie_core_clk_clk),                                            //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                       //                     reset.reset
		.uav_address              (sgdma_m_read_translator_avalon_universal_master_0_address),            // avalon_universal_master_0.address
		.uav_burstcount           (sgdma_m_read_translator_avalon_universal_master_0_burstcount),         //                          .burstcount
		.uav_read                 (sgdma_m_read_translator_avalon_universal_master_0_read),               //                          .read
		.uav_write                (sgdma_m_read_translator_avalon_universal_master_0_write),              //                          .write
		.uav_waitrequest          (sgdma_m_read_translator_avalon_universal_master_0_waitrequest),        //                          .waitrequest
		.uav_readdatavalid        (sgdma_m_read_translator_avalon_universal_master_0_readdatavalid),      //                          .readdatavalid
		.uav_byteenable           (sgdma_m_read_translator_avalon_universal_master_0_byteenable),         //                          .byteenable
		.uav_readdata             (sgdma_m_read_translator_avalon_universal_master_0_readdata),           //                          .readdata
		.uav_writedata            (sgdma_m_read_translator_avalon_universal_master_0_writedata),          //                          .writedata
		.uav_lock                 (sgdma_m_read_translator_avalon_universal_master_0_lock),               //                          .lock
		.uav_debugaccess          (sgdma_m_read_translator_avalon_universal_master_0_debugaccess),        //                          .debugaccess
		.av_address               (sgdma_m_read_address),                                                 //      avalon_anti_master_0.address
		.av_waitrequest           (sgdma_m_read_waitrequest),                                             //                          .waitrequest
		.av_burstcount            (sgdma_m_read_burstcount),                                              //                          .burstcount
		.av_read                  (sgdma_m_read_read),                                                    //                          .read
		.av_readdata              (sgdma_m_read_readdata),                                                //                          .readdata
		.av_readdatavalid         (sgdma_m_read_readdatavalid),                                           //                          .readdatavalid
		.av_byteenable            (8'b11111111),                                                          //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                 //               (terminated)
		.av_begintransfer         (1'b0),                                                                 //               (terminated)
		.av_chipselect            (1'b0),                                                                 //               (terminated)
		.av_write                 (1'b0),                                                                 //               (terminated)
		.av_writedata             (64'b0000000000000000000000000000000000000000000000000000000000000000), //               (terminated)
		.av_lock                  (1'b0),                                                                 //               (terminated)
		.av_debugaccess           (1'b0),                                                                 //               (terminated)
		.uav_clken                (),                                                                     //               (terminated)
		.av_clken                 (1'b1),                                                                 //               (terminated)
		.uav_response             (2'b00),                                                                //               (terminated)
		.av_response              (),                                                                     //               (terminated)
		.uav_writeresponserequest (),                                                                     //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                 //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                 //               (terminated)
		.av_writeresponsevalid    ()                                                                      //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (64),
		.AV_BURSTCOUNT_W             (8),
		.AV_BYTEENABLE_W             (8),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (11),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (8),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (1),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_m_write_translator (
		.clk                      (pcie_ip_pcie_core_clk_clk),                                        //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                   //                     reset.reset
		.uav_address              (sgdma_m_write_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (sgdma_m_write_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (sgdma_m_write_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (sgdma_m_write_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (sgdma_m_write_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (sgdma_m_write_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (sgdma_m_write_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (sgdma_m_write_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (sgdma_m_write_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (sgdma_m_write_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (sgdma_m_write_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (sgdma_m_write_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (sgdma_m_write_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (sgdma_m_write_burstcount),                                         //                          .burstcount
		.av_byteenable            (sgdma_m_write_byteenable),                                         //                          .byteenable
		.av_write                 (sgdma_m_write_write),                                              //                          .write
		.av_writedata             (sgdma_m_write_writedata),                                          //                          .writedata
		.av_beginbursttransfer    (1'b0),                                                             //               (terminated)
		.av_begintransfer         (1'b0),                                                             //               (terminated)
		.av_chipselect            (1'b0),                                                             //               (terminated)
		.av_read                  (1'b0),                                                             //               (terminated)
		.av_readdata              (),                                                                 //               (terminated)
		.av_readdatavalid         (),                                                                 //               (terminated)
		.av_lock                  (1'b0),                                                             //               (terminated)
		.av_debugaccess           (1'b0),                                                             //               (terminated)
		.uav_clken                (),                                                                 //               (terminated)
		.av_clken                 (1'b1),                                                             //               (terminated)
		.uav_response             (2'b00),                                                            //               (terminated)
		.av_response              (),                                                                 //               (terminated)
		.uav_writeresponserequest (),                                                                 //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                             //               (terminated)
		.av_writeresponserequest  (1'b0),                                                             //               (terminated)
		.av_writeresponsevalid    ()                                                                  //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (31),
		.AV_DATA_W                      (64),
		.UAV_DATA_W                     (64),
		.AV_BURSTCOUNT_W                (7),
		.AV_BYTEENABLE_W                (8),
		.UAV_BYTEENABLE_W               (8),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (10),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (8),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pcie_ip_txs_translator (
		.clk                      (pcie_ip_pcie_core_clk_clk),                                              //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                     //                    reset.reset
		.uav_address              (pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pcie_ip_txs_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (pcie_ip_txs_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (pcie_ip_txs_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (pcie_ip_txs_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (pcie_ip_txs_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount            (pcie_ip_txs_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable            (pcie_ip_txs_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (pcie_ip_txs_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (pcie_ip_txs_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (pcie_ip_txs_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (24),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_s1_translator (
		.clk                      (clk_clk),                                                             //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                  //                    reset.reset
		.uav_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sdram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sdram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (sdram_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (sdram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sdram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (sdram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (sdram_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (sdram_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (sdram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (64),
		.AV_BURSTCOUNT_W             (7),
		.AV_BYTEENABLE_W             (8),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (10),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (8),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (1),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) pcie_ip_bar1_0_translator (
		.clk                      (pcie_ip_pcie_core_clk_clk),                                         //                       clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                //                     reset.reset
		.uav_address              (pcie_ip_bar1_0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (pcie_ip_bar1_0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (pcie_ip_bar1_0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (pcie_ip_bar1_0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (pcie_ip_bar1_0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (pcie_ip_bar1_0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (pcie_ip_bar1_0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (pcie_ip_bar1_0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (pcie_ip_bar1_0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (pcie_ip_bar1_0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (pcie_ip_bar1_0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (pcie_ip_bar1_0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (pcie_ip_bar1_0_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (pcie_ip_bar1_0_burstcount),                                         //                          .burstcount
		.av_byteenable            (pcie_ip_bar1_0_byteenable),                                         //                          .byteenable
		.av_read                  (pcie_ip_bar1_0_read),                                               //                          .read
		.av_readdata              (pcie_ip_bar1_0_readdata),                                           //                          .readdata
		.av_readdatavalid         (pcie_ip_bar1_0_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (pcie_ip_bar1_0_write),                                              //                          .write
		.av_writedata             (pcie_ip_bar1_0_writedata),                                          //                          .writedata
		.av_beginbursttransfer    (1'b0),                                                              //               (terminated)
		.av_begintransfer         (1'b0),                                                              //               (terminated)
		.av_chipselect            (1'b0),                                                              //               (terminated)
		.av_lock                  (1'b0),                                                              //               (terminated)
		.av_debugaccess           (1'b0),                                                              //               (terminated)
		.uav_clken                (),                                                                  //               (terminated)
		.av_clken                 (1'b1),                                                              //               (terminated)
		.uav_response             (2'b00),                                                             //               (terminated)
		.av_response              (),                                                                  //               (terminated)
		.uav_writeresponserequest (),                                                                  //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                              //               (terminated)
		.av_writeresponserequest  (1'b0),                                                              //               (terminated)
		.av_writeresponsevalid    ()                                                                   //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (5),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) custom_slave_block_0_avalon_slave_translator (
		.clk                      (clk_clk),                                                                                      //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                                           //                    reset.reset
		.uav_address              (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (custom_slave_block_0_avalon_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (custom_slave_block_0_avalon_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (custom_slave_block_0_avalon_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (custom_slave_block_0_avalon_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (custom_slave_block_0_avalon_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (custom_slave_block_0_avalon_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                                             //              (terminated)
		.av_burstcount            (),                                                                                             //              (terminated)
		.av_byteenable            (),                                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                                             //              (terminated)
		.av_lock                  (),                                                                                             //              (terminated)
		.av_clken                 (),                                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                                         //              (terminated)
		.av_debugaccess           (),                                                                                             //              (terminated)
		.av_outputenable          (),                                                                                             //              (terminated)
		.uav_response             (),                                                                                             //              (terminated)
		.av_response              (2'b00),                                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                          //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (135),
		.PKT_PROTECTION_L          (133),
		.PKT_BEGIN_BURST           (128),
		.PKT_BURSTWRAP_H           (120),
		.PKT_BURSTWRAP_L           (120),
		.PKT_BURST_SIZE_H          (123),
		.PKT_BURST_SIZE_L          (121),
		.PKT_BURST_TYPE_H          (125),
		.PKT_BURST_TYPE_L          (124),
		.PKT_BYTE_CNT_H            (119),
		.PKT_BYTE_CNT_L            (110),
		.PKT_ADDR_H                (103),
		.PKT_ADDR_L                (72),
		.PKT_TRANS_COMPRESSED_READ (104),
		.PKT_TRANS_POSTED          (105),
		.PKT_TRANS_WRITE           (106),
		.PKT_TRANS_READ            (107),
		.PKT_TRANS_LOCK            (108),
		.PKT_TRANS_EXCLUSIVE       (109),
		.PKT_DATA_H                (63),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64),
		.PKT_SRC_ID_H              (130),
		.PKT_SRC_ID_L              (130),
		.PKT_DEST_ID_H             (131),
		.PKT_DEST_ID_L             (131),
		.PKT_THREAD_ID_H           (132),
		.PKT_THREAD_ID_L           (132),
		.PKT_CACHE_H               (139),
		.PKT_CACHE_L               (136),
		.PKT_DATA_SIDEBAND_H       (127),
		.PKT_DATA_SIDEBAND_L       (127),
		.PKT_QOS_H                 (129),
		.PKT_QOS_L                 (129),
		.PKT_ADDR_SIDEBAND_H       (126),
		.PKT_ADDR_SIDEBAND_L       (126),
		.PKT_RESPONSE_STATUS_H     (141),
		.PKT_RESPONSE_STATUS_L     (140),
		.ST_DATA_W                 (142),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (10),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pcie_ip_bar2_translator_avalon_universal_master_0_agent (
		.clk                     (pcie_ip_pcie_core_clk_clk),                                                //       clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                       // clk_reset.reset
		.av_address              (pcie_ip_bar2_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (pcie_ip_bar2_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (pcie_ip_bar2_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (pcie_ip_bar2_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (pcie_ip_bar2_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (pcie_ip_bar2_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (pcie_ip_bar2_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (pcie_ip_bar2_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (pcie_ip_bar2_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (pcie_ip_bar2_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (pcie_ip_bar2_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (pcie_ip_bar2_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (pcie_ip_bar2_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (pcie_ip_bar2_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (pcie_ip_bar2_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (pcie_ip_bar2_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_rsp_src_valid),                                                    //        rp.valid
		.rp_data                 (limiter_rsp_src_data),                                                     //          .data
		.rp_channel              (limiter_rsp_src_channel),                                                  //          .channel
		.rp_startofpacket        (limiter_rsp_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket          (limiter_rsp_src_endofpacket),                                              //          .endofpacket
		.rp_ready                (limiter_rsp_src_ready),                                                    //          .ready
		.av_response             (),                                                                         // (terminated)
		.av_writeresponserequest (1'b0),                                                                     // (terminated)
		.av_writeresponsevalid   ()                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (95),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (84),
		.PKT_BYTE_CNT_H            (83),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (99),
		.PKT_PROTECTION_L          (97),
		.PKT_RESPONSE_STATUS_H     (105),
		.PKT_RESPONSE_STATUS_L     (104),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (106),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sgdma_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (pcie_ip_pcie_core_clk_clk),                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (sgdma_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sgdma_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sgdma_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sgdma_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sgdma_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sgdma_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sgdma_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sgdma_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sgdma_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sgdma_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sgdma_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sgdma_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sgdma_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sgdma_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sgdma_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sgdma_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                    //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                    //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                     //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                              //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                  //                .channel
		.rf_sink_ready           (sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sgdma_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sgdma_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sgdma_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sgdma_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sgdma_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sgdma_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (107),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pcie_ip_pcie_core_clk_clk),                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sgdma_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sgdma_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (95),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (84),
		.PKT_BYTE_CNT_H            (83),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (99),
		.PKT_PROTECTION_L          (97),
		.PKT_RESPONSE_STATUS_H     (105),
		.PKT_RESPONSE_STATUS_L     (104),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (106),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pcie_ip_cra_translator_avalon_universal_slave_0_agent (
		.clk                     (pcie_ip_pcie_core_clk_clk),                                                        //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pcie_ip_cra_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                                  //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                                  //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                   //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                            //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                                //                .channel
		.rf_sink_ready           (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (107),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pcie_ip_pcie_core_clk_clk),                                                        //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                               // clk_reset.reset
		.in_data           (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_BEGIN_BURST           (93),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (85),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.PKT_BURST_TYPE_H          (90),
		.PKT_BURST_TYPE_L          (89),
		.PKT_BYTE_CNT_H            (84),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (96),
		.PKT_SRC_ID_L              (95),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (97),
		.PKT_THREAD_ID_H           (99),
		.PKT_THREAD_ID_L           (99),
		.PKT_CACHE_H               (106),
		.PKT_CACHE_L               (103),
		.PKT_DATA_SIDEBAND_H       (92),
		.PKT_DATA_SIDEBAND_L       (92),
		.PKT_QOS_H                 (94),
		.PKT_QOS_L                 (94),
		.PKT_ADDR_SIDEBAND_H       (91),
		.PKT_ADDR_SIDEBAND_L       (91),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.ST_DATA_W                 (109),
		.ST_CHANNEL_W              (4),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (0),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sgdma_descriptor_read_translator_avalon_universal_master_0_agent (
		.clk                     (pcie_ip_pcie_core_clk_clk),                                                         //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.av_address              (sgdma_descriptor_read_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (sgdma_descriptor_read_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (sgdma_descriptor_read_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (sgdma_descriptor_read_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (sgdma_descriptor_read_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (sgdma_descriptor_read_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (sgdma_descriptor_read_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (sgdma_descriptor_read_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (sgdma_descriptor_read_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (sgdma_descriptor_read_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (sgdma_descriptor_read_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (width_adapter_008_src_valid),                                                       //        rp.valid
		.rp_data                 (width_adapter_008_src_data),                                                        //          .data
		.rp_channel              (width_adapter_008_src_channel),                                                     //          .channel
		.rp_startofpacket        (width_adapter_008_src_startofpacket),                                               //          .startofpacket
		.rp_endofpacket          (width_adapter_008_src_endofpacket),                                                 //          .endofpacket
		.rp_ready                (width_adapter_008_src_ready),                                                       //          .ready
		.av_response             (),                                                                                  // (terminated)
		.av_writeresponserequest (1'b0),                                                                              // (terminated)
		.av_writeresponsevalid   ()                                                                                   // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_BEGIN_BURST           (93),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (85),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.PKT_BURST_TYPE_H          (90),
		.PKT_BURST_TYPE_L          (89),
		.PKT_BYTE_CNT_H            (84),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (96),
		.PKT_SRC_ID_L              (95),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (97),
		.PKT_THREAD_ID_H           (99),
		.PKT_THREAD_ID_L           (99),
		.PKT_CACHE_H               (106),
		.PKT_CACHE_L               (103),
		.PKT_DATA_SIDEBAND_H       (92),
		.PKT_DATA_SIDEBAND_L       (92),
		.PKT_QOS_H                 (94),
		.PKT_QOS_L                 (94),
		.PKT_ADDR_SIDEBAND_H       (91),
		.PKT_ADDR_SIDEBAND_L       (91),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.ST_DATA_W                 (109),
		.ST_CHANNEL_W              (4),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (1),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sgdma_descriptor_write_translator_avalon_universal_master_0_agent (
		.clk                     (pcie_ip_pcie_core_clk_clk),                                                          //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.av_address              (sgdma_descriptor_write_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (sgdma_descriptor_write_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (sgdma_descriptor_write_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (sgdma_descriptor_write_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (sgdma_descriptor_write_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (sgdma_descriptor_write_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (sgdma_descriptor_write_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (sgdma_descriptor_write_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (sgdma_descriptor_write_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (sgdma_descriptor_write_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (sgdma_descriptor_write_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (width_adapter_009_src_valid),                                                        //        rp.valid
		.rp_data                 (width_adapter_009_src_data),                                                         //          .data
		.rp_channel              (width_adapter_009_src_channel),                                                      //          .channel
		.rp_startofpacket        (width_adapter_009_src_startofpacket),                                                //          .startofpacket
		.rp_endofpacket          (width_adapter_009_src_endofpacket),                                                  //          .endofpacket
		.rp_ready                (width_adapter_009_src_ready),                                                        //          .ready
		.av_response             (),                                                                                   // (terminated)
		.av_writeresponserequest (1'b0),                                                                               // (terminated)
		.av_writeresponsevalid   ()                                                                                    // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (138),
		.PKT_PROTECTION_L          (136),
		.PKT_BEGIN_BURST           (129),
		.PKT_BURSTWRAP_H           (121),
		.PKT_BURSTWRAP_L           (121),
		.PKT_BURST_SIZE_H          (124),
		.PKT_BURST_SIZE_L          (122),
		.PKT_BURST_TYPE_H          (126),
		.PKT_BURST_TYPE_L          (125),
		.PKT_BYTE_CNT_H            (120),
		.PKT_BYTE_CNT_L            (110),
		.PKT_ADDR_H                (103),
		.PKT_ADDR_L                (72),
		.PKT_TRANS_COMPRESSED_READ (104),
		.PKT_TRANS_POSTED          (105),
		.PKT_TRANS_WRITE           (106),
		.PKT_TRANS_READ            (107),
		.PKT_TRANS_LOCK            (108),
		.PKT_TRANS_EXCLUSIVE       (109),
		.PKT_DATA_H                (63),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64),
		.PKT_SRC_ID_H              (132),
		.PKT_SRC_ID_L              (131),
		.PKT_DEST_ID_H             (134),
		.PKT_DEST_ID_L             (133),
		.PKT_THREAD_ID_H           (135),
		.PKT_THREAD_ID_L           (135),
		.PKT_CACHE_H               (142),
		.PKT_CACHE_L               (139),
		.PKT_DATA_SIDEBAND_H       (128),
		.PKT_DATA_SIDEBAND_L       (128),
		.PKT_QOS_H                 (130),
		.PKT_QOS_L                 (130),
		.PKT_ADDR_SIDEBAND_H       (127),
		.PKT_ADDR_SIDEBAND_L       (127),
		.PKT_RESPONSE_STATUS_H     (144),
		.PKT_RESPONSE_STATUS_L     (143),
		.ST_DATA_W                 (145),
		.ST_CHANNEL_W              (4),
		.AV_BURSTCOUNT_W           (7),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sgdma_m_read_translator_avalon_universal_master_0_agent (
		.clk                     (pcie_ip_pcie_core_clk_clk),                                                //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.av_address              (sgdma_m_read_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (sgdma_m_read_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (sgdma_m_read_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (sgdma_m_read_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (sgdma_m_read_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (sgdma_m_read_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (sgdma_m_read_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (sgdma_m_read_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (sgdma_m_read_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (sgdma_m_read_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (sgdma_m_read_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (sgdma_m_read_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (sgdma_m_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (sgdma_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (sgdma_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (sgdma_m_read_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_001_rsp_src_valid),                                                //        rp.valid
		.rp_data                 (limiter_001_rsp_src_data),                                                 //          .data
		.rp_channel              (limiter_001_rsp_src_channel),                                              //          .channel
		.rp_startofpacket        (limiter_001_rsp_src_startofpacket),                                        //          .startofpacket
		.rp_endofpacket          (limiter_001_rsp_src_endofpacket),                                          //          .endofpacket
		.rp_ready                (limiter_001_rsp_src_ready),                                                //          .ready
		.av_response             (),                                                                         // (terminated)
		.av_writeresponserequest (1'b0),                                                                     // (terminated)
		.av_writeresponsevalid   ()                                                                          // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (138),
		.PKT_PROTECTION_L          (136),
		.PKT_BEGIN_BURST           (129),
		.PKT_BURSTWRAP_H           (121),
		.PKT_BURSTWRAP_L           (121),
		.PKT_BURST_SIZE_H          (124),
		.PKT_BURST_SIZE_L          (122),
		.PKT_BURST_TYPE_H          (126),
		.PKT_BURST_TYPE_L          (125),
		.PKT_BYTE_CNT_H            (120),
		.PKT_BYTE_CNT_L            (110),
		.PKT_ADDR_H                (103),
		.PKT_ADDR_L                (72),
		.PKT_TRANS_COMPRESSED_READ (104),
		.PKT_TRANS_POSTED          (105),
		.PKT_TRANS_WRITE           (106),
		.PKT_TRANS_READ            (107),
		.PKT_TRANS_LOCK            (108),
		.PKT_TRANS_EXCLUSIVE       (109),
		.PKT_DATA_H                (63),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64),
		.PKT_SRC_ID_H              (132),
		.PKT_SRC_ID_L              (131),
		.PKT_DEST_ID_H             (134),
		.PKT_DEST_ID_L             (133),
		.PKT_THREAD_ID_H           (135),
		.PKT_THREAD_ID_L           (135),
		.PKT_CACHE_H               (142),
		.PKT_CACHE_L               (139),
		.PKT_DATA_SIDEBAND_H       (128),
		.PKT_DATA_SIDEBAND_L       (128),
		.PKT_QOS_H                 (130),
		.PKT_QOS_L                 (130),
		.PKT_ADDR_SIDEBAND_H       (127),
		.PKT_ADDR_SIDEBAND_L       (127),
		.PKT_RESPONSE_STATUS_H     (144),
		.PKT_RESPONSE_STATUS_L     (143),
		.ST_DATA_W                 (145),
		.ST_CHANNEL_W              (4),
		.AV_BURSTCOUNT_W           (11),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (3),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sgdma_m_write_translator_avalon_universal_master_0_agent (
		.clk                     (pcie_ip_pcie_core_clk_clk),                                                 //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                            // clk_reset.reset
		.av_address              (sgdma_m_write_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (sgdma_m_write_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (sgdma_m_write_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (sgdma_m_write_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (sgdma_m_write_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (sgdma_m_write_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (sgdma_m_write_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (sgdma_m_write_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (sgdma_m_write_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (sgdma_m_write_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (sgdma_m_write_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (sgdma_m_write_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (sgdma_m_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (sgdma_m_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (sgdma_m_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (sgdma_m_write_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_004_src_valid),                                                //        rp.valid
		.rp_data                 (rsp_xbar_mux_004_src_data),                                                 //          .data
		.rp_channel              (rsp_xbar_mux_004_src_channel),                                              //          .channel
		.rp_startofpacket        (rsp_xbar_mux_004_src_startofpacket),                                        //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_004_src_endofpacket),                                          //          .endofpacket
		.rp_ready                (rsp_xbar_mux_004_src_ready),                                                //          .ready
		.av_response             (),                                                                          // (terminated)
		.av_writeresponserequest (1'b0),                                                                      // (terminated)
		.av_writeresponsevalid   ()                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (63),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (129),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64),
		.PKT_ADDR_H                (103),
		.PKT_ADDR_L                (72),
		.PKT_TRANS_COMPRESSED_READ (104),
		.PKT_TRANS_POSTED          (105),
		.PKT_TRANS_WRITE           (106),
		.PKT_TRANS_READ            (107),
		.PKT_TRANS_LOCK            (108),
		.PKT_SRC_ID_H              (132),
		.PKT_SRC_ID_L              (131),
		.PKT_DEST_ID_H             (134),
		.PKT_DEST_ID_L             (133),
		.PKT_BURSTWRAP_H           (121),
		.PKT_BURSTWRAP_L           (121),
		.PKT_BYTE_CNT_H            (120),
		.PKT_BYTE_CNT_L            (110),
		.PKT_PROTECTION_H          (138),
		.PKT_PROTECTION_L          (136),
		.PKT_RESPONSE_STATUS_H     (144),
		.PKT_RESPONSE_STATUS_L     (143),
		.PKT_BURST_SIZE_H          (124),
		.PKT_BURST_SIZE_L          (122),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (145),
		.AVS_BURSTCOUNT_W          (10),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pcie_ip_txs_translator_avalon_universal_slave_0_agent (
		.clk                     (pcie_ip_pcie_core_clk_clk),                                                        //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pcie_ip_txs_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_002_source0_ready),                                                  //              cp.ready
		.cp_valid                (burst_adapter_002_source0_valid),                                                  //                .valid
		.cp_data                 (burst_adapter_002_source0_data),                                                   //                .data
		.cp_startofpacket        (burst_adapter_002_source0_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (burst_adapter_002_source0_endofpacket),                                            //                .endofpacket
		.cp_channel              (burst_adapter_002_source0_channel),                                                //                .channel
		.rf_sink_ready           (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (146),
		.FIFO_DEPTH          (9),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pcie_ip_pcie_core_clk_clk),                                                        //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                               // clk_reset.reset
		.in_data           (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (93),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (96),
		.PKT_SRC_ID_L              (95),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (97),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (85),
		.PKT_BYTE_CNT_H            (84),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_003_source0_ready),                                               //              cp.ready
		.cp_valid                (burst_adapter_003_source0_valid),                                               //                .valid
		.cp_data                 (burst_adapter_003_source0_data),                                                //                .data
		.cp_startofpacket        (burst_adapter_003_source0_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (burst_adapter_003_source0_endofpacket),                                         //                .endofpacket
		.cp_channel              (burst_adapter_003_source0_channel),                                             //                .channel
		.rf_sink_ready           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                       //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                   // (terminated)
		.csr_read          (1'b0),                                                                    // (terminated)
		.csr_write         (1'b0),                                                                    // (terminated)
		.csr_readdata      (),                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                    // (terminated)
		.almost_full_data  (),                                                                        // (terminated)
		.almost_empty_data (),                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                    // (terminated)
		.out_startofpacket (),                                                                        // (terminated)
		.out_endofpacket   (),                                                                        // (terminated)
		.in_empty          (1'b0),                                                                    // (terminated)
		.out_empty         (),                                                                        // (terminated)
		.in_error          (1'b0),                                                                    // (terminated)
		.out_error         (),                                                                        // (terminated)
		.in_channel        (1'b0),                                                                    // (terminated)
		.out_channel       ()                                                                         // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (135),
		.PKT_PROTECTION_L          (133),
		.PKT_BEGIN_BURST           (128),
		.PKT_BURSTWRAP_H           (120),
		.PKT_BURSTWRAP_L           (120),
		.PKT_BURST_SIZE_H          (123),
		.PKT_BURST_SIZE_L          (121),
		.PKT_BURST_TYPE_H          (125),
		.PKT_BURST_TYPE_L          (124),
		.PKT_BYTE_CNT_H            (119),
		.PKT_BYTE_CNT_L            (110),
		.PKT_ADDR_H                (103),
		.PKT_ADDR_L                (72),
		.PKT_TRANS_COMPRESSED_READ (104),
		.PKT_TRANS_POSTED          (105),
		.PKT_TRANS_WRITE           (106),
		.PKT_TRANS_READ            (107),
		.PKT_TRANS_LOCK            (108),
		.PKT_TRANS_EXCLUSIVE       (109),
		.PKT_DATA_H                (63),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64),
		.PKT_SRC_ID_H              (130),
		.PKT_SRC_ID_L              (130),
		.PKT_DEST_ID_H             (131),
		.PKT_DEST_ID_L             (131),
		.PKT_THREAD_ID_H           (132),
		.PKT_THREAD_ID_L           (132),
		.PKT_CACHE_H               (139),
		.PKT_CACHE_L               (136),
		.PKT_DATA_SIDEBAND_H       (127),
		.PKT_DATA_SIDEBAND_L       (127),
		.PKT_QOS_H                 (129),
		.PKT_QOS_L                 (129),
		.PKT_ADDR_SIDEBAND_H       (126),
		.PKT_ADDR_SIDEBAND_L       (126),
		.PKT_RESPONSE_STATUS_H     (141),
		.PKT_RESPONSE_STATUS_L     (140),
		.ST_DATA_W                 (142),
		.ST_CHANNEL_W              (1),
		.AV_BURSTCOUNT_W           (10),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pcie_ip_bar1_0_translator_avalon_universal_master_0_agent (
		.clk                     (pcie_ip_pcie_core_clk_clk),                                                  //       clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                         // clk_reset.reset
		.av_address              (pcie_ip_bar1_0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (pcie_ip_bar1_0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (pcie_ip_bar1_0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (pcie_ip_bar1_0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (pcie_ip_bar1_0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (pcie_ip_bar1_0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (pcie_ip_bar1_0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (pcie_ip_bar1_0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (pcie_ip_bar1_0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (pcie_ip_bar1_0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (pcie_ip_bar1_0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (pcie_ip_bar1_0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (pcie_ip_bar1_0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (pcie_ip_bar1_0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (pcie_ip_bar1_0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (pcie_ip_bar1_0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (crosser_001_out_valid),                                                      //        rp.valid
		.rp_data                 (crosser_001_out_data),                                                       //          .data
		.rp_channel              (crosser_001_out_channel),                                                    //          .channel
		.rp_startofpacket        (crosser_001_out_startofpacket),                                              //          .startofpacket
		.rp_endofpacket          (crosser_001_out_endofpacket),                                                //          .endofpacket
		.rp_ready                (crosser_001_out_ready),                                                      //          .ready
		.av_response             (),                                                                           // (terminated)
		.av_writeresponserequest (1'b0),                                                                       // (terminated)
		.av_writeresponsevalid   ()                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (95),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (84),
		.PKT_BYTE_CNT_H            (83),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (99),
		.PKT_PROTECTION_L          (97),
		.PKT_RESPONSE_STATUS_H     (105),
		.PKT_RESPONSE_STATUS_L     (104),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (1),
		.ST_DATA_W                 (106),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                                //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_004_source0_ready),                                                                        //              cp.ready
		.cp_valid                (burst_adapter_004_source0_valid),                                                                        //                .valid
		.cp_data                 (burst_adapter_004_source0_data),                                                                         //                .data
		.cp_startofpacket        (burst_adapter_004_source0_startofpacket),                                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_004_source0_endofpacket),                                                                  //                .endofpacket
		.cp_channel              (burst_adapter_004_source0_channel),                                                                      //                .channel
		.rf_sink_ready           (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (107),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                                //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                                   // (terminated)
		.csr_readdata      (),                                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                   // (terminated)
		.almost_full_data  (),                                                                                                       // (terminated)
		.almost_empty_data (),                                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                                   // (terminated)
		.out_empty         (),                                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                                   // (terminated)
		.out_error         (),                                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                                   // (terminated)
		.out_channel       ()                                                                                                        // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                                          //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_startofpacket  (1'b0),                                                                                             // (terminated)
		.in_endofpacket    (1'b0),                                                                                             // (terminated)
		.out_startofpacket (),                                                                                                 // (terminated)
		.out_endofpacket   (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	amm_master_qsys_with_pcie_addr_router addr_router (
		.sink_ready         (pcie_ip_bar2_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (pcie_ip_bar2_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (pcie_ip_bar2_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (pcie_ip_bar2_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pcie_ip_bar2_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pcie_ip_pcie_core_clk_clk),                                                //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                    //       src.ready
		.src_valid          (addr_router_src_valid),                                                    //          .valid
		.src_data           (addr_router_src_data),                                                     //          .data
		.src_channel        (addr_router_src_channel),                                                  //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                               //          .endofpacket
	);

	amm_master_qsys_with_pcie_id_router id_router (
		.sink_ready         (sgdma_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sgdma_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sgdma_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sgdma_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pcie_ip_pcie_core_clk_clk),                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                  //       src.ready
		.src_valid          (id_router_src_valid),                                                  //          .valid
		.src_data           (id_router_src_data),                                                   //          .data
		.src_channel        (id_router_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                             //          .endofpacket
	);

	amm_master_qsys_with_pcie_id_router id_router_001 (
		.sink_ready         (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pcie_ip_cra_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pcie_ip_pcie_core_clk_clk),                                              //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                //       src.ready
		.src_valid          (id_router_001_src_valid),                                                //          .valid
		.src_data           (id_router_001_src_data),                                                 //          .data
		.src_channel        (id_router_001_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                           //          .endofpacket
	);

	amm_master_qsys_with_pcie_addr_router_001 addr_router_001 (
		.sink_ready         (sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pcie_ip_pcie_core_clk_clk),                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                         //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                         //          .valid
		.src_data           (addr_router_001_src_data),                                                          //          .data
		.src_channel        (addr_router_001_src_channel),                                                       //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                    //          .endofpacket
	);

	amm_master_qsys_with_pcie_addr_router_001 addr_router_002 (
		.sink_ready         (sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pcie_ip_pcie_core_clk_clk),                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                          //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                          //          .valid
		.src_data           (addr_router_002_src_data),                                                           //          .data
		.src_channel        (addr_router_002_src_channel),                                                        //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                     //          .endofpacket
	);

	amm_master_qsys_with_pcie_addr_router_003 addr_router_003 (
		.sink_ready         (sgdma_m_read_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_m_read_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_m_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pcie_ip_pcie_core_clk_clk),                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                //          .valid
		.src_data           (addr_router_003_src_data),                                                 //          .data
		.src_channel        (addr_router_003_src_channel),                                              //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                           //          .endofpacket
	);

	amm_master_qsys_with_pcie_addr_router_003 addr_router_004 (
		.sink_ready         (sgdma_m_write_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_m_write_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_m_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_m_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_m_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pcie_ip_pcie_core_clk_clk),                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (addr_router_004_src_ready),                                                 //       src.ready
		.src_valid          (addr_router_004_src_valid),                                                 //          .valid
		.src_data           (addr_router_004_src_data),                                                  //          .data
		.src_channel        (addr_router_004_src_channel),                                               //          .channel
		.src_startofpacket  (addr_router_004_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (addr_router_004_src_endofpacket)                                            //          .endofpacket
	);

	amm_master_qsys_with_pcie_id_router_002 id_router_002 (
		.sink_ready         (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pcie_ip_txs_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pcie_ip_pcie_core_clk_clk),                                              //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                //       src.ready
		.src_valid          (id_router_002_src_valid),                                                //          .valid
		.src_data           (id_router_002_src_data),                                                 //          .data
		.src_channel        (id_router_002_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                           //          .endofpacket
	);

	amm_master_qsys_with_pcie_id_router_003 id_router_003 (
		.sink_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                             //       src.ready
		.src_valid          (id_router_003_src_valid),                                             //          .valid
		.src_data           (id_router_003_src_data),                                              //          .data
		.src_channel        (id_router_003_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                        //          .endofpacket
	);

	amm_master_qsys_with_pcie_addr_router_005 addr_router_005 (
		.sink_ready         (pcie_ip_bar1_0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (pcie_ip_bar1_0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (pcie_ip_bar1_0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (pcie_ip_bar1_0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pcie_ip_bar1_0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pcie_ip_pcie_core_clk_clk),                                                  //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (addr_router_005_src_ready),                                                  //       src.ready
		.src_valid          (addr_router_005_src_valid),                                                  //          .valid
		.src_data           (addr_router_005_src_data),                                                   //          .data
		.src_channel        (addr_router_005_src_channel),                                                //          .channel
		.src_startofpacket  (addr_router_005_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (addr_router_005_src_endofpacket)                                             //          .endofpacket
	);

	amm_master_qsys_with_pcie_id_router_004 id_router_004 (
		.sink_ready         (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (custom_slave_block_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                      //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                                      //       src.ready
		.src_valid          (id_router_004_src_valid),                                                                      //          .valid
		.src_data           (id_router_004_src_data),                                                                       //          .data
		.src_channel        (id_router_004_src_channel),                                                                    //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                              //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                                 //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (131),
		.PKT_DEST_ID_L             (131),
		.PKT_TRANS_POSTED          (105),
		.PKT_TRANS_WRITE           (106),
		.MAX_OUTSTANDING_RESPONSES (3),
		.PIPELINED                 (0),
		.ST_DATA_W                 (142),
		.ST_CHANNEL_W              (2),
		.VALID_WIDTH               (2),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (119),
		.PKT_BYTE_CNT_L            (110),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64)
	) limiter (
		.clk                    (pcie_ip_pcie_core_clk_clk),          //       clk.clk
		.reset                  (rst_controller_003_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),              //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),              //          .valid
		.cmd_sink_data          (addr_router_src_data),               //          .data
		.cmd_sink_channel       (addr_router_src_channel),            //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),      //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),        //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),              //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),               //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),            //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),      //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),        //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),             //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),             //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),           //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),              //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket),     //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),       //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),              //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),              //          .valid
		.rsp_src_data           (limiter_rsp_src_data),               //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),            //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),      //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),        //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)              // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (134),
		.PKT_DEST_ID_L             (133),
		.PKT_TRANS_POSTED          (105),
		.PKT_TRANS_WRITE           (106),
		.MAX_OUTSTANDING_RESPONSES (13),
		.PIPELINED                 (0),
		.ST_DATA_W                 (145),
		.ST_CHANNEL_W              (4),
		.VALID_WIDTH               (4),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (120),
		.PKT_BYTE_CNT_L            (110),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64)
	) limiter_001 (
		.clk                    (pcie_ip_pcie_core_clk_clk),          //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_003_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_003_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_003_src_data),           //          .data
		.cmd_sink_channel       (addr_router_003_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_003_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_003_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_003_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_003_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_003_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_003_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_003_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_003_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (92),
		.PKT_BYTE_CNT_H            (83),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.PKT_BURST_TYPE_H          (89),
		.PKT_BURST_TYPE_L          (88),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (84),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (106),
		.ST_CHANNEL_W              (2),
		.OUT_BYTE_CNT_H            (76),
		.OUT_BURSTWRAP_H           (84),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (1),
		.BURSTWRAP_CONST_VALUE     (1)
	) burst_adapter (
		.clk                   (pcie_ip_pcie_core_clk_clk),           //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_src_data),              //          .data
		.sink0_channel         (width_adapter_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),             //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (92),
		.PKT_BYTE_CNT_H            (83),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.PKT_BURST_TYPE_H          (89),
		.PKT_BURST_TYPE_L          (88),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (84),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (106),
		.ST_CHANNEL_W              (2),
		.OUT_BYTE_CNT_H            (76),
		.OUT_BURSTWRAP_H           (84),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (1),
		.BURSTWRAP_CONST_VALUE     (1)
	) burst_adapter_001 (
		.clk                   (pcie_ip_pcie_core_clk_clk),               //       cr0.clk
		.reset                 (rst_controller_003_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (width_adapter_002_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_002_src_data),              //          .data
		.sink0_channel         (width_adapter_002_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_002_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_002_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_002_src_ready),             //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (103),
		.PKT_ADDR_L                (72),
		.PKT_BEGIN_BURST           (129),
		.PKT_BYTE_CNT_H            (120),
		.PKT_BYTE_CNT_L            (110),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64),
		.PKT_BURST_SIZE_H          (124),
		.PKT_BURST_SIZE_L          (122),
		.PKT_BURST_TYPE_H          (126),
		.PKT_BURST_TYPE_L          (125),
		.PKT_BURSTWRAP_H           (121),
		.PKT_BURSTWRAP_L           (121),
		.PKT_TRANS_COMPRESSED_READ (104),
		.PKT_TRANS_WRITE           (106),
		.PKT_TRANS_READ            (107),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (145),
		.ST_CHANNEL_W              (4),
		.OUT_BYTE_CNT_H            (119),
		.OUT_BURSTWRAP_H           (121),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (1),
		.BURSTWRAP_CONST_VALUE     (1)
	) burst_adapter_002 (
		.clk                   (pcie_ip_pcie_core_clk_clk),               //       cr0.clk
		.reset                 (rst_controller_003_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_002_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_002_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_002_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_002_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_002_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_002_src_ready),              //          .ready
		.source0_valid         (burst_adapter_002_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_002_source0_data),          //          .data
		.source0_channel       (burst_adapter_002_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_002_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_002_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_002_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (93),
		.PKT_BYTE_CNT_H            (84),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (88),
		.PKT_BURST_SIZE_L          (86),
		.PKT_BURST_TYPE_H          (90),
		.PKT_BURST_TYPE_L          (89),
		.PKT_BURSTWRAP_H           (85),
		.PKT_BURSTWRAP_L           (85),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (109),
		.ST_CHANNEL_W              (4),
		.OUT_BYTE_CNT_H            (76),
		.OUT_BURSTWRAP_H           (85),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (1),
		.BURSTWRAP_CONST_VALUE     (1)
	) burst_adapter_003 (
		.clk                   (clk_clk),                                 //       cr0.clk
		.reset                 (rst_controller_001_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_003_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_003_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_003_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_003_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_003_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_003_src_ready),              //          .ready
		.source0_valid         (burst_adapter_003_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_003_source0_data),          //          .data
		.source0_channel       (burst_adapter_003_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_003_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_003_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_003_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (92),
		.PKT_BYTE_CNT_H            (83),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.PKT_BURST_TYPE_H          (89),
		.PKT_BURST_TYPE_L          (88),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (84),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (106),
		.ST_CHANNEL_W              (1),
		.OUT_BYTE_CNT_H            (76),
		.OUT_BURSTWRAP_H           (84),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (1),
		.BURSTWRAP_CONST_VALUE     (1)
	) burst_adapter_004 (
		.clk                   (clk_clk),                                 //       cr0.clk
		.reset                 (rst_controller_002_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (width_adapter_012_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_012_src_data),              //          .data
		.sink0_channel         (width_adapter_012_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_012_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_012_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_012_src_ready),             //          .ready
		.source0_valid         (burst_adapter_004_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_004_source0_data),          //          .data
		.source0_channel       (burst_adapter_004_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_004_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_004_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_004_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.reset_in1  (~pcie_ip_pcie_core_reset_reset), // reset_in1.reset
		.clk        (pcie_ip_pcie_core_clk_clk),      //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.reset_in1  (~pcie_ip_pcie_core_reset_reset),     // reset_in1.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_002 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_003 (
		.reset_in0  (~pcie_ip_pcie_core_reset_reset),     // reset_in0.reset
		.clk        (pcie_ip_pcie_core_clk_clk),          //       clk.clk
		.reset_out  (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	amm_master_qsys_with_pcie_cmd_xbar_demux cmd_xbar_demux (
		.clk                (pcie_ip_pcie_core_clk_clk),          //        clk.clk
		.reset              (rst_controller_003_reset_out_reset), //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),              //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),            //           .channel
		.sink_data          (limiter_cmd_src_data),               //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),             // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),          //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),          //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),           //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),        //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),    //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),          //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),          //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),           //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),        //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket)     //           .endofpacket
	);

	amm_master_qsys_with_pcie_rsp_xbar_demux rsp_xbar_demux (
		.clk                (pcie_ip_pcie_core_clk_clk),           //       clk.clk
		.reset              (rst_controller_reset_out_reset),      // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),         //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),       //          .channel
		.sink_data          (width_adapter_001_src_data),          //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket), //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),   //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),         //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),           //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),           //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),            //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),         //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket),   //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket)      //          .endofpacket
	);

	amm_master_qsys_with_pcie_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (pcie_ip_pcie_core_clk_clk),             //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (width_adapter_003_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_003_src_channel),         //          .channel
		.sink_data          (width_adapter_003_src_data),            //          .data
		.sink_startofpacket (width_adapter_003_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_003_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_003_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	amm_master_qsys_with_pcie_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (pcie_ip_pcie_core_clk_clk),             //       clk.clk
		.reset               (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	amm_master_qsys_with_pcie_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (pcie_ip_pcie_core_clk_clk),             //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	amm_master_qsys_with_pcie_cmd_xbar_demux_001 cmd_xbar_demux_002 (
		.clk                (pcie_ip_pcie_core_clk_clk),             //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_002_src_ready),             //      sink.ready
		.sink_channel       (addr_router_002_src_channel),           //          .channel
		.sink_data          (addr_router_002_src_data),              //          .data
		.sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_002_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	amm_master_qsys_with_pcie_cmd_xbar_demux_003 cmd_xbar_demux_003 (
		.clk                (pcie_ip_pcie_core_clk_clk),             //        clk.clk
		.reset              (rst_controller_reset_out_reset),        //  clk_reset.reset
		.sink_ready         (limiter_001_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_001_cmd_src_channel),           //           .channel
		.sink_data          (limiter_001_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_001_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_001_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_001_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_003_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_003_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_003_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_003_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_003_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_003_src1_endofpacket)    //           .endofpacket
	);

	amm_master_qsys_with_pcie_cmd_xbar_demux_004 cmd_xbar_demux_004 (
		.clk                (pcie_ip_pcie_core_clk_clk),             //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_004_src_ready),             //      sink.ready
		.sink_channel       (addr_router_004_src_channel),           //          .channel
		.sink_data          (addr_router_004_src_data),              //          .data
		.sink_startofpacket (addr_router_004_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_004_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_004_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_004_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_004_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_004_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_004_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_004_src1_endofpacket)    //          .endofpacket
	);

	amm_master_qsys_with_pcie_cmd_xbar_mux_002 cmd_xbar_mux_002 (
		.clk                 (pcie_ip_pcie_core_clk_clk),             //       clk.clk
		.reset               (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (width_adapter_004_src_ready),           //     sink0.ready
		.sink0_valid         (width_adapter_004_src_valid),           //          .valid
		.sink0_channel       (width_adapter_004_src_channel),         //          .channel
		.sink0_data          (width_adapter_004_src_data),            //          .data
		.sink0_startofpacket (width_adapter_004_src_startofpacket),   //          .startofpacket
		.sink0_endofpacket   (width_adapter_004_src_endofpacket),     //          .endofpacket
		.sink1_ready         (width_adapter_005_src_ready),           //     sink1.ready
		.sink1_valid         (width_adapter_005_src_valid),           //          .valid
		.sink1_channel       (width_adapter_005_src_channel),         //          .channel
		.sink1_data          (width_adapter_005_src_data),            //          .data
		.sink1_startofpacket (width_adapter_005_src_startofpacket),   //          .startofpacket
		.sink1_endofpacket   (width_adapter_005_src_endofpacket),     //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_003_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_004_src0_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_004_src0_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_004_src0_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_004_src0_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	amm_master_qsys_with_pcie_cmd_xbar_mux_003 cmd_xbar_mux_003 (
		.clk                 (clk_clk),                            //       clk.clk
		.reset               (rst_controller_001_reset_out_reset), // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),         //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),         //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),          //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),       //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket), //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),   //          .endofpacket
		.sink0_ready         (crosser_002_out_ready),              //     sink0.ready
		.sink0_valid         (crosser_002_out_valid),              //          .valid
		.sink0_channel       (crosser_002_out_channel),            //          .channel
		.sink0_data          (crosser_002_out_data),               //          .data
		.sink0_startofpacket (crosser_002_out_startofpacket),      //          .startofpacket
		.sink0_endofpacket   (crosser_002_out_endofpacket),        //          .endofpacket
		.sink1_ready         (crosser_003_out_ready),              //     sink1.ready
		.sink1_valid         (crosser_003_out_valid),              //          .valid
		.sink1_channel       (crosser_003_out_channel),            //          .channel
		.sink1_data          (crosser_003_out_data),               //          .data
		.sink1_startofpacket (crosser_003_out_startofpacket),      //          .startofpacket
		.sink1_endofpacket   (crosser_003_out_endofpacket)         //          .endofpacket
	);

	amm_master_qsys_with_pcie_rsp_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (pcie_ip_pcie_core_clk_clk),             //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_002_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_002_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_002_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_002_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_002_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_002_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_002_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_002_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_002_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_002_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_002_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_002_src3_endofpacket)    //          .endofpacket
	);

	amm_master_qsys_with_pcie_rsp_xbar_demux_003 rsp_xbar_demux_003 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	amm_master_qsys_with_pcie_rsp_xbar_mux_003 rsp_xbar_mux_003 (
		.clk                 (pcie_ip_pcie_core_clk_clk),             //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_003_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_003_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_002_src2_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_002_src2_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_002_src2_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_002_src2_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_002_src2_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_002_src2_endofpacket),   //          .endofpacket
		.sink1_ready         (crosser_004_out_ready),                 //     sink1.ready
		.sink1_valid         (crosser_004_out_valid),                 //          .valid
		.sink1_channel       (crosser_004_out_channel),               //          .channel
		.sink1_data          (crosser_004_out_data),                  //          .data
		.sink1_startofpacket (crosser_004_out_startofpacket),         //          .startofpacket
		.sink1_endofpacket   (crosser_004_out_endofpacket)            //          .endofpacket
	);

	amm_master_qsys_with_pcie_rsp_xbar_mux_003 rsp_xbar_mux_004 (
		.clk                 (pcie_ip_pcie_core_clk_clk),             //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_004_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_004_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_004_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_004_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_004_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_004_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_002_src3_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_002_src3_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_002_src3_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_002_src3_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_002_src3_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_002_src3_endofpacket),   //          .endofpacket
		.sink1_ready         (crosser_005_out_ready),                 //     sink1.ready
		.sink1_valid         (crosser_005_out_valid),                 //          .valid
		.sink1_channel       (crosser_005_out_channel),               //          .channel
		.sink1_data          (crosser_005_out_data),                  //          .data
		.sink1_startofpacket (crosser_005_out_startofpacket),         //          .startofpacket
		.sink1_endofpacket   (crosser_005_out_endofpacket)            //          .endofpacket
	);

	amm_master_qsys_with_pcie_cmd_xbar_demux_005 cmd_xbar_demux_005 (
		.clk                (pcie_ip_pcie_core_clk_clk),             //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_005_src_ready),             //      sink.ready
		.sink_channel       (addr_router_005_src_channel),           //          .channel
		.sink_data          (addr_router_005_src_data),              //          .data
		.sink_startofpacket (addr_router_005_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_005_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_005_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	amm_master_qsys_with_pcie_cmd_xbar_demux_005 rsp_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (width_adapter_013_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_013_src_channel),         //          .channel
		.sink_data          (width_adapter_013_src_data),            //          .data
		.sink_startofpacket (width_adapter_013_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_013_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_013_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (103),
		.IN_PKT_ADDR_L                 (72),
		.IN_PKT_DATA_H                 (63),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (71),
		.IN_PKT_BYTEEN_L               (64),
		.IN_PKT_BYTE_CNT_H             (119),
		.IN_PKT_BYTE_CNT_L             (110),
		.IN_PKT_TRANS_COMPRESSED_READ  (104),
		.IN_PKT_BURSTWRAP_H            (120),
		.IN_PKT_BURSTWRAP_L            (120),
		.IN_PKT_BURST_SIZE_H           (123),
		.IN_PKT_BURST_SIZE_L           (121),
		.IN_PKT_RESPONSE_STATUS_H      (141),
		.IN_PKT_RESPONSE_STATUS_L      (140),
		.IN_PKT_TRANS_EXCLUSIVE        (109),
		.IN_PKT_BURST_TYPE_H           (125),
		.IN_PKT_BURST_TYPE_L           (124),
		.IN_ST_DATA_W                  (142),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (83),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (87),
		.OUT_PKT_BURST_SIZE_L          (85),
		.OUT_PKT_RESPONSE_STATUS_H     (105),
		.OUT_PKT_RESPONSE_STATUS_L     (104),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (89),
		.OUT_PKT_BURST_TYPE_L          (88),
		.OUT_ST_DATA_W                 (106),
		.ST_CHANNEL_W                  (2),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter (
		.clk                  (pcie_ip_pcie_core_clk_clk),         //       clk.clk
		.reset                (rst_controller_reset_out_reset),    // clk_reset.reset
		.in_valid             (cmd_xbar_demux_src0_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_src0_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_src0_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_src0_ready),         //          .ready
		.in_data              (cmd_xbar_demux_src0_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_src_data),            //          .data
		.out_channel          (width_adapter_src_channel),         //          .channel
		.out_valid            (width_adapter_src_valid),           //          .valid
		.out_ready            (width_adapter_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                             // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (83),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (84),
		.IN_PKT_BURSTWRAP_L            (84),
		.IN_PKT_BURST_SIZE_H           (87),
		.IN_PKT_BURST_SIZE_L           (85),
		.IN_PKT_RESPONSE_STATUS_H      (105),
		.IN_PKT_RESPONSE_STATUS_L      (104),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (89),
		.IN_PKT_BURST_TYPE_L           (88),
		.IN_ST_DATA_W                  (106),
		.OUT_PKT_ADDR_H                (103),
		.OUT_PKT_ADDR_L                (72),
		.OUT_PKT_DATA_H                (63),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (71),
		.OUT_PKT_BYTEEN_L              (64),
		.OUT_PKT_BYTE_CNT_H            (119),
		.OUT_PKT_BYTE_CNT_L            (110),
		.OUT_PKT_TRANS_COMPRESSED_READ (104),
		.OUT_PKT_BURST_SIZE_H          (123),
		.OUT_PKT_BURST_SIZE_L          (121),
		.OUT_PKT_RESPONSE_STATUS_H     (141),
		.OUT_PKT_RESPONSE_STATUS_L     (140),
		.OUT_PKT_TRANS_EXCLUSIVE       (109),
		.OUT_PKT_BURST_TYPE_H          (125),
		.OUT_PKT_BURST_TYPE_L          (124),
		.OUT_ST_DATA_W                 (142),
		.ST_CHANNEL_W                  (2),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (1)
	) width_adapter_001 (
		.clk                  (pcie_ip_pcie_core_clk_clk),           //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_src_valid),                 //      sink.valid
		.in_channel           (id_router_src_channel),               //          .channel
		.in_startofpacket     (id_router_src_startofpacket),         //          .startofpacket
		.in_endofpacket       (id_router_src_endofpacket),           //          .endofpacket
		.in_ready             (id_router_src_ready),                 //          .ready
		.in_data              (id_router_src_data),                  //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (103),
		.IN_PKT_ADDR_L                 (72),
		.IN_PKT_DATA_H                 (63),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (71),
		.IN_PKT_BYTEEN_L               (64),
		.IN_PKT_BYTE_CNT_H             (119),
		.IN_PKT_BYTE_CNT_L             (110),
		.IN_PKT_TRANS_COMPRESSED_READ  (104),
		.IN_PKT_BURSTWRAP_H            (120),
		.IN_PKT_BURSTWRAP_L            (120),
		.IN_PKT_BURST_SIZE_H           (123),
		.IN_PKT_BURST_SIZE_L           (121),
		.IN_PKT_RESPONSE_STATUS_H      (141),
		.IN_PKT_RESPONSE_STATUS_L      (140),
		.IN_PKT_TRANS_EXCLUSIVE        (109),
		.IN_PKT_BURST_TYPE_H           (125),
		.IN_PKT_BURST_TYPE_L           (124),
		.IN_ST_DATA_W                  (142),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (83),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (87),
		.OUT_PKT_BURST_SIZE_L          (85),
		.OUT_PKT_RESPONSE_STATUS_H     (105),
		.OUT_PKT_RESPONSE_STATUS_L     (104),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (89),
		.OUT_PKT_BURST_TYPE_L          (88),
		.OUT_ST_DATA_W                 (106),
		.ST_CHANNEL_W                  (2),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_002 (
		.clk                  (pcie_ip_pcie_core_clk_clk),           //       clk.clk
		.reset                (rst_controller_003_reset_out_reset),  // clk_reset.reset
		.in_valid             (cmd_xbar_demux_src1_valid),           //      sink.valid
		.in_channel           (cmd_xbar_demux_src1_channel),         //          .channel
		.in_startofpacket     (cmd_xbar_demux_src1_startofpacket),   //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_src1_endofpacket),     //          .endofpacket
		.in_ready             (cmd_xbar_demux_src1_ready),           //          .ready
		.in_data              (cmd_xbar_demux_src1_data),            //          .data
		.out_endofpacket      (width_adapter_002_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_002_src_data),          //          .data
		.out_channel          (width_adapter_002_src_channel),       //          .channel
		.out_valid            (width_adapter_002_src_valid),         //          .valid
		.out_ready            (width_adapter_002_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_002_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (83),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (84),
		.IN_PKT_BURSTWRAP_L            (84),
		.IN_PKT_BURST_SIZE_H           (87),
		.IN_PKT_BURST_SIZE_L           (85),
		.IN_PKT_RESPONSE_STATUS_H      (105),
		.IN_PKT_RESPONSE_STATUS_L      (104),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (89),
		.IN_PKT_BURST_TYPE_L           (88),
		.IN_ST_DATA_W                  (106),
		.OUT_PKT_ADDR_H                (103),
		.OUT_PKT_ADDR_L                (72),
		.OUT_PKT_DATA_H                (63),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (71),
		.OUT_PKT_BYTEEN_L              (64),
		.OUT_PKT_BYTE_CNT_H            (119),
		.OUT_PKT_BYTE_CNT_L            (110),
		.OUT_PKT_TRANS_COMPRESSED_READ (104),
		.OUT_PKT_BURST_SIZE_H          (123),
		.OUT_PKT_BURST_SIZE_L          (121),
		.OUT_PKT_RESPONSE_STATUS_H     (141),
		.OUT_PKT_RESPONSE_STATUS_L     (140),
		.OUT_PKT_TRANS_EXCLUSIVE       (109),
		.OUT_PKT_BURST_TYPE_H          (125),
		.OUT_PKT_BURST_TYPE_L          (124),
		.OUT_ST_DATA_W                 (142),
		.ST_CHANNEL_W                  (2),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (1)
	) width_adapter_003 (
		.clk                  (pcie_ip_pcie_core_clk_clk),           //       clk.clk
		.reset                (rst_controller_003_reset_out_reset),  // clk_reset.reset
		.in_valid             (id_router_001_src_valid),             //      sink.valid
		.in_channel           (id_router_001_src_channel),           //          .channel
		.in_startofpacket     (id_router_001_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_001_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_001_src_ready),             //          .ready
		.in_data              (id_router_001_src_data),              //          .data
		.out_endofpacket      (width_adapter_003_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_003_src_data),          //          .data
		.out_channel          (width_adapter_003_src_channel),       //          .channel
		.out_valid            (width_adapter_003_src_valid),         //          .valid
		.out_ready            (width_adapter_003_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_003_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (84),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (85),
		.IN_PKT_BURSTWRAP_L            (85),
		.IN_PKT_BURST_SIZE_H           (88),
		.IN_PKT_BURST_SIZE_L           (86),
		.IN_PKT_RESPONSE_STATUS_H      (108),
		.IN_PKT_RESPONSE_STATUS_L      (107),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (90),
		.IN_PKT_BURST_TYPE_L           (89),
		.IN_ST_DATA_W                  (109),
		.OUT_PKT_ADDR_H                (103),
		.OUT_PKT_ADDR_L                (72),
		.OUT_PKT_DATA_H                (63),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (71),
		.OUT_PKT_BYTEEN_L              (64),
		.OUT_PKT_BYTE_CNT_H            (120),
		.OUT_PKT_BYTE_CNT_L            (110),
		.OUT_PKT_TRANS_COMPRESSED_READ (104),
		.OUT_PKT_BURST_SIZE_H          (124),
		.OUT_PKT_BURST_SIZE_L          (122),
		.OUT_PKT_RESPONSE_STATUS_H     (144),
		.OUT_PKT_RESPONSE_STATUS_L     (143),
		.OUT_PKT_TRANS_EXCLUSIVE       (109),
		.OUT_PKT_BURST_TYPE_H          (126),
		.OUT_PKT_BURST_TYPE_L          (125),
		.OUT_ST_DATA_W                 (145),
		.ST_CHANNEL_W                  (4),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_004 (
		.clk                  (pcie_ip_pcie_core_clk_clk),             //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src0_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src0_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src0_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src0_data),          //          .data
		.out_endofpacket      (width_adapter_004_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_004_src_data),            //          .data
		.out_channel          (width_adapter_004_src_channel),         //          .channel
		.out_valid            (width_adapter_004_src_valid),           //          .valid
		.out_ready            (width_adapter_004_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_004_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (84),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (85),
		.IN_PKT_BURSTWRAP_L            (85),
		.IN_PKT_BURST_SIZE_H           (88),
		.IN_PKT_BURST_SIZE_L           (86),
		.IN_PKT_RESPONSE_STATUS_H      (108),
		.IN_PKT_RESPONSE_STATUS_L      (107),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (90),
		.IN_PKT_BURST_TYPE_L           (89),
		.IN_ST_DATA_W                  (109),
		.OUT_PKT_ADDR_H                (103),
		.OUT_PKT_ADDR_L                (72),
		.OUT_PKT_DATA_H                (63),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (71),
		.OUT_PKT_BYTEEN_L              (64),
		.OUT_PKT_BYTE_CNT_H            (120),
		.OUT_PKT_BYTE_CNT_L            (110),
		.OUT_PKT_TRANS_COMPRESSED_READ (104),
		.OUT_PKT_BURST_SIZE_H          (124),
		.OUT_PKT_BURST_SIZE_L          (122),
		.OUT_PKT_RESPONSE_STATUS_H     (144),
		.OUT_PKT_RESPONSE_STATUS_L     (143),
		.OUT_PKT_TRANS_EXCLUSIVE       (109),
		.OUT_PKT_BURST_TYPE_H          (126),
		.OUT_PKT_BURST_TYPE_L          (125),
		.OUT_ST_DATA_W                 (145),
		.ST_CHANNEL_W                  (4),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_005 (
		.clk                  (pcie_ip_pcie_core_clk_clk),             //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_002_src0_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_002_src0_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_002_src0_ready),         //          .ready
		.in_data              (cmd_xbar_demux_002_src0_data),          //          .data
		.out_endofpacket      (width_adapter_005_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_005_src_data),            //          .data
		.out_channel          (width_adapter_005_src_channel),         //          .channel
		.out_valid            (width_adapter_005_src_valid),           //          .valid
		.out_ready            (width_adapter_005_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_005_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (103),
		.IN_PKT_ADDR_L                 (72),
		.IN_PKT_DATA_H                 (63),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (71),
		.IN_PKT_BYTEEN_L               (64),
		.IN_PKT_BYTE_CNT_H             (120),
		.IN_PKT_BYTE_CNT_L             (110),
		.IN_PKT_TRANS_COMPRESSED_READ  (104),
		.IN_PKT_BURSTWRAP_H            (121),
		.IN_PKT_BURSTWRAP_L            (121),
		.IN_PKT_BURST_SIZE_H           (124),
		.IN_PKT_BURST_SIZE_L           (122),
		.IN_PKT_RESPONSE_STATUS_H      (144),
		.IN_PKT_RESPONSE_STATUS_L      (143),
		.IN_PKT_TRANS_EXCLUSIVE        (109),
		.IN_PKT_BURST_TYPE_H           (126),
		.IN_PKT_BURST_TYPE_L           (125),
		.IN_ST_DATA_W                  (145),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (84),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (88),
		.OUT_PKT_BURST_SIZE_L          (86),
		.OUT_PKT_RESPONSE_STATUS_H     (108),
		.OUT_PKT_RESPONSE_STATUS_L     (107),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (90),
		.OUT_PKT_BURST_TYPE_L          (89),
		.OUT_ST_DATA_W                 (109),
		.ST_CHANNEL_W                  (4),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_006 (
		.clk                  (pcie_ip_pcie_core_clk_clk),             //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_003_src1_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_003_src1_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_003_src1_ready),         //          .ready
		.in_data              (cmd_xbar_demux_003_src1_data),          //          .data
		.out_endofpacket      (width_adapter_006_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_006_src_data),            //          .data
		.out_channel          (width_adapter_006_src_channel),         //          .channel
		.out_valid            (width_adapter_006_src_valid),           //          .valid
		.out_ready            (width_adapter_006_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_006_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (103),
		.IN_PKT_ADDR_L                 (72),
		.IN_PKT_DATA_H                 (63),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (71),
		.IN_PKT_BYTEEN_L               (64),
		.IN_PKT_BYTE_CNT_H             (120),
		.IN_PKT_BYTE_CNT_L             (110),
		.IN_PKT_TRANS_COMPRESSED_READ  (104),
		.IN_PKT_BURSTWRAP_H            (121),
		.IN_PKT_BURSTWRAP_L            (121),
		.IN_PKT_BURST_SIZE_H           (124),
		.IN_PKT_BURST_SIZE_L           (122),
		.IN_PKT_RESPONSE_STATUS_H      (144),
		.IN_PKT_RESPONSE_STATUS_L      (143),
		.IN_PKT_TRANS_EXCLUSIVE        (109),
		.IN_PKT_BURST_TYPE_H           (126),
		.IN_PKT_BURST_TYPE_L           (125),
		.IN_ST_DATA_W                  (145),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (84),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (88),
		.OUT_PKT_BURST_SIZE_L          (86),
		.OUT_PKT_RESPONSE_STATUS_H     (108),
		.OUT_PKT_RESPONSE_STATUS_L     (107),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (90),
		.OUT_PKT_BURST_TYPE_L          (89),
		.OUT_ST_DATA_W                 (109),
		.ST_CHANNEL_W                  (4),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_007 (
		.clk                  (pcie_ip_pcie_core_clk_clk),             //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_004_src1_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_004_src1_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_004_src1_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_004_src1_ready),         //          .ready
		.in_data              (cmd_xbar_demux_004_src1_data),          //          .data
		.out_endofpacket      (width_adapter_007_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_007_src_data),            //          .data
		.out_channel          (width_adapter_007_src_channel),         //          .channel
		.out_valid            (width_adapter_007_src_valid),           //          .valid
		.out_ready            (width_adapter_007_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_007_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (103),
		.IN_PKT_ADDR_L                 (72),
		.IN_PKT_DATA_H                 (63),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (71),
		.IN_PKT_BYTEEN_L               (64),
		.IN_PKT_BYTE_CNT_H             (120),
		.IN_PKT_BYTE_CNT_L             (110),
		.IN_PKT_TRANS_COMPRESSED_READ  (104),
		.IN_PKT_BURSTWRAP_H            (121),
		.IN_PKT_BURSTWRAP_L            (121),
		.IN_PKT_BURST_SIZE_H           (124),
		.IN_PKT_BURST_SIZE_L           (122),
		.IN_PKT_RESPONSE_STATUS_H      (144),
		.IN_PKT_RESPONSE_STATUS_L      (143),
		.IN_PKT_TRANS_EXCLUSIVE        (109),
		.IN_PKT_BURST_TYPE_H           (126),
		.IN_PKT_BURST_TYPE_L           (125),
		.IN_ST_DATA_W                  (145),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (84),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (88),
		.OUT_PKT_BURST_SIZE_L          (86),
		.OUT_PKT_RESPONSE_STATUS_H     (108),
		.OUT_PKT_RESPONSE_STATUS_L     (107),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (90),
		.OUT_PKT_BURST_TYPE_L          (89),
		.OUT_ST_DATA_W                 (109),
		.ST_CHANNEL_W                  (4),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_008 (
		.clk                  (pcie_ip_pcie_core_clk_clk),             //       clk.clk
		.reset                (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.in_valid             (rsp_xbar_demux_002_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_002_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_002_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_002_src0_data),          //          .data
		.out_endofpacket      (width_adapter_008_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_008_src_data),            //          .data
		.out_channel          (width_adapter_008_src_channel),         //          .channel
		.out_valid            (width_adapter_008_src_valid),           //          .valid
		.out_ready            (width_adapter_008_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_008_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (103),
		.IN_PKT_ADDR_L                 (72),
		.IN_PKT_DATA_H                 (63),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (71),
		.IN_PKT_BYTEEN_L               (64),
		.IN_PKT_BYTE_CNT_H             (120),
		.IN_PKT_BYTE_CNT_L             (110),
		.IN_PKT_TRANS_COMPRESSED_READ  (104),
		.IN_PKT_BURSTWRAP_H            (121),
		.IN_PKT_BURSTWRAP_L            (121),
		.IN_PKT_BURST_SIZE_H           (124),
		.IN_PKT_BURST_SIZE_L           (122),
		.IN_PKT_RESPONSE_STATUS_H      (144),
		.IN_PKT_RESPONSE_STATUS_L      (143),
		.IN_PKT_TRANS_EXCLUSIVE        (109),
		.IN_PKT_BURST_TYPE_H           (126),
		.IN_PKT_BURST_TYPE_L           (125),
		.IN_ST_DATA_W                  (145),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (84),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (88),
		.OUT_PKT_BURST_SIZE_L          (86),
		.OUT_PKT_RESPONSE_STATUS_H     (108),
		.OUT_PKT_RESPONSE_STATUS_L     (107),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (90),
		.OUT_PKT_BURST_TYPE_L          (89),
		.OUT_ST_DATA_W                 (109),
		.ST_CHANNEL_W                  (4),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_009 (
		.clk                  (pcie_ip_pcie_core_clk_clk),             //       clk.clk
		.reset                (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.in_valid             (rsp_xbar_demux_002_src1_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_002_src1_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_002_src1_ready),         //          .ready
		.in_data              (rsp_xbar_demux_002_src1_data),          //          .data
		.out_endofpacket      (width_adapter_009_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_009_src_data),            //          .data
		.out_channel          (width_adapter_009_src_channel),         //          .channel
		.out_valid            (width_adapter_009_src_valid),           //          .valid
		.out_ready            (width_adapter_009_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_009_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (84),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (85),
		.IN_PKT_BURSTWRAP_L            (85),
		.IN_PKT_BURST_SIZE_H           (88),
		.IN_PKT_BURST_SIZE_L           (86),
		.IN_PKT_RESPONSE_STATUS_H      (108),
		.IN_PKT_RESPONSE_STATUS_L      (107),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (90),
		.IN_PKT_BURST_TYPE_L           (89),
		.IN_ST_DATA_W                  (109),
		.OUT_PKT_ADDR_H                (103),
		.OUT_PKT_ADDR_L                (72),
		.OUT_PKT_DATA_H                (63),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (71),
		.OUT_PKT_BYTEEN_L              (64),
		.OUT_PKT_BYTE_CNT_H            (120),
		.OUT_PKT_BYTE_CNT_L            (110),
		.OUT_PKT_TRANS_COMPRESSED_READ (104),
		.OUT_PKT_BURST_SIZE_H          (124),
		.OUT_PKT_BURST_SIZE_L          (122),
		.OUT_PKT_RESPONSE_STATUS_H     (144),
		.OUT_PKT_RESPONSE_STATUS_L     (143),
		.OUT_PKT_TRANS_EXCLUSIVE       (109),
		.OUT_PKT_BURST_TYPE_H          (126),
		.OUT_PKT_BURST_TYPE_L          (125),
		.OUT_ST_DATA_W                 (145),
		.ST_CHANNEL_W                  (4),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (1)
	) width_adapter_010 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.in_valid             (rsp_xbar_demux_003_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_003_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_003_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_003_src0_data),          //          .data
		.out_endofpacket      (width_adapter_010_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_010_src_data),            //          .data
		.out_channel          (width_adapter_010_src_channel),         //          .channel
		.out_valid            (width_adapter_010_src_valid),           //          .valid
		.out_ready            (width_adapter_010_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_010_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (84),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (85),
		.IN_PKT_BURSTWRAP_L            (85),
		.IN_PKT_BURST_SIZE_H           (88),
		.IN_PKT_BURST_SIZE_L           (86),
		.IN_PKT_RESPONSE_STATUS_H      (108),
		.IN_PKT_RESPONSE_STATUS_L      (107),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (90),
		.IN_PKT_BURST_TYPE_L           (89),
		.IN_ST_DATA_W                  (109),
		.OUT_PKT_ADDR_H                (103),
		.OUT_PKT_ADDR_L                (72),
		.OUT_PKT_DATA_H                (63),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (71),
		.OUT_PKT_BYTEEN_L              (64),
		.OUT_PKT_BYTE_CNT_H            (120),
		.OUT_PKT_BYTE_CNT_L            (110),
		.OUT_PKT_TRANS_COMPRESSED_READ (104),
		.OUT_PKT_BURST_SIZE_H          (124),
		.OUT_PKT_BURST_SIZE_L          (122),
		.OUT_PKT_RESPONSE_STATUS_H     (144),
		.OUT_PKT_RESPONSE_STATUS_L     (143),
		.OUT_PKT_TRANS_EXCLUSIVE       (109),
		.OUT_PKT_BURST_TYPE_H          (126),
		.OUT_PKT_BURST_TYPE_L          (125),
		.OUT_ST_DATA_W                 (145),
		.ST_CHANNEL_W                  (4),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (1)
	) width_adapter_011 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.in_valid             (rsp_xbar_demux_003_src1_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_003_src1_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_003_src1_ready),         //          .ready
		.in_data              (rsp_xbar_demux_003_src1_data),          //          .data
		.out_endofpacket      (width_adapter_011_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_011_src_data),            //          .data
		.out_channel          (width_adapter_011_src_channel),         //          .channel
		.out_valid            (width_adapter_011_src_valid),           //          .valid
		.out_ready            (width_adapter_011_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_011_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (103),
		.IN_PKT_ADDR_L                 (72),
		.IN_PKT_DATA_H                 (63),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (71),
		.IN_PKT_BYTEEN_L               (64),
		.IN_PKT_BYTE_CNT_H             (119),
		.IN_PKT_BYTE_CNT_L             (110),
		.IN_PKT_TRANS_COMPRESSED_READ  (104),
		.IN_PKT_BURSTWRAP_H            (120),
		.IN_PKT_BURSTWRAP_L            (120),
		.IN_PKT_BURST_SIZE_H           (123),
		.IN_PKT_BURST_SIZE_L           (121),
		.IN_PKT_RESPONSE_STATUS_H      (141),
		.IN_PKT_RESPONSE_STATUS_L      (140),
		.IN_PKT_TRANS_EXCLUSIVE        (109),
		.IN_PKT_BURST_TYPE_H           (125),
		.IN_PKT_BURST_TYPE_L           (124),
		.IN_ST_DATA_W                  (142),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (83),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (87),
		.OUT_PKT_BURST_SIZE_L          (85),
		.OUT_PKT_RESPONSE_STATUS_H     (105),
		.OUT_PKT_RESPONSE_STATUS_L     (104),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (89),
		.OUT_PKT_BURST_TYPE_L          (88),
		.OUT_ST_DATA_W                 (106),
		.ST_CHANNEL_W                  (1),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_012 (
		.clk                  (clk_clk),                             //       clk.clk
		.reset                (rst_controller_002_reset_out_reset),  // clk_reset.reset
		.in_valid             (crosser_out_valid),                   //      sink.valid
		.in_channel           (crosser_out_channel),                 //          .channel
		.in_startofpacket     (crosser_out_startofpacket),           //          .startofpacket
		.in_endofpacket       (crosser_out_endofpacket),             //          .endofpacket
		.in_ready             (crosser_out_ready),                   //          .ready
		.in_data              (crosser_out_data),                    //          .data
		.out_endofpacket      (width_adapter_012_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_012_src_data),          //          .data
		.out_channel          (width_adapter_012_src_channel),       //          .channel
		.out_valid            (width_adapter_012_src_valid),         //          .valid
		.out_ready            (width_adapter_012_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_012_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (83),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (84),
		.IN_PKT_BURSTWRAP_L            (84),
		.IN_PKT_BURST_SIZE_H           (87),
		.IN_PKT_BURST_SIZE_L           (85),
		.IN_PKT_RESPONSE_STATUS_H      (105),
		.IN_PKT_RESPONSE_STATUS_L      (104),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (89),
		.IN_PKT_BURST_TYPE_L           (88),
		.IN_ST_DATA_W                  (106),
		.OUT_PKT_ADDR_H                (103),
		.OUT_PKT_ADDR_L                (72),
		.OUT_PKT_DATA_H                (63),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (71),
		.OUT_PKT_BYTEEN_L              (64),
		.OUT_PKT_BYTE_CNT_H            (119),
		.OUT_PKT_BYTE_CNT_L            (110),
		.OUT_PKT_TRANS_COMPRESSED_READ (104),
		.OUT_PKT_BURST_SIZE_H          (123),
		.OUT_PKT_BURST_SIZE_L          (121),
		.OUT_PKT_RESPONSE_STATUS_H     (141),
		.OUT_PKT_RESPONSE_STATUS_L     (140),
		.OUT_PKT_TRANS_EXCLUSIVE       (109),
		.OUT_PKT_BURST_TYPE_H          (125),
		.OUT_PKT_BURST_TYPE_L          (124),
		.OUT_ST_DATA_W                 (142),
		.ST_CHANNEL_W                  (1),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (1)
	) width_adapter_013 (
		.clk                  (clk_clk),                             //       clk.clk
		.reset                (rst_controller_002_reset_out_reset),  // clk_reset.reset
		.in_valid             (id_router_004_src_valid),             //      sink.valid
		.in_channel           (id_router_004_src_channel),           //          .channel
		.in_startofpacket     (id_router_004_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_004_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_004_src_ready),             //          .ready
		.in_data              (id_router_004_src_data),              //          .data
		.out_endofpacket      (width_adapter_013_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_013_src_data),          //          .data
		.out_channel          (width_adapter_013_src_channel),       //          .channel
		.out_valid            (width_adapter_013_src_valid),         //          .valid
		.out_ready            (width_adapter_013_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_013_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (142),
		.BITS_PER_SYMBOL     (142),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (1),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (pcie_ip_pcie_core_clk_clk),             //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_002_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_005_src0_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_005_src0_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_005_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_005_src0_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_005_src0_channel),       //              .channel
		.in_data           (cmd_xbar_demux_005_src0_data),          //              .data
		.out_ready         (crosser_out_ready),                     //           out.ready
		.out_valid         (crosser_out_valid),                     //              .valid
		.out_startofpacket (crosser_out_startofpacket),             //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),               //              .endofpacket
		.out_channel       (crosser_out_channel),                   //              .channel
		.out_data          (crosser_out_data),                      //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (142),
		.BITS_PER_SYMBOL     (142),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (1),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_002_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (pcie_ip_pcie_core_clk_clk),             //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_004_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_004_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_004_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_004_src0_data),          //              .data
		.out_ready         (crosser_001_out_ready),                 //           out.ready
		.out_valid         (crosser_001_out_valid),                 //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_001_out_channel),               //              .channel
		.out_data          (crosser_001_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (109),
		.BITS_PER_SYMBOL     (109),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (4),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_002 (
		.in_clk            (pcie_ip_pcie_core_clk_clk),           //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),      //  in_clk_reset.reset
		.out_clk           (clk_clk),                             //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),  // out_clk_reset.reset
		.in_ready          (width_adapter_006_src_ready),         //            in.ready
		.in_valid          (width_adapter_006_src_valid),         //              .valid
		.in_startofpacket  (width_adapter_006_src_startofpacket), //              .startofpacket
		.in_endofpacket    (width_adapter_006_src_endofpacket),   //              .endofpacket
		.in_channel        (width_adapter_006_src_channel),       //              .channel
		.in_data           (width_adapter_006_src_data),          //              .data
		.out_ready         (crosser_002_out_ready),               //           out.ready
		.out_valid         (crosser_002_out_valid),               //              .valid
		.out_startofpacket (crosser_002_out_startofpacket),       //              .startofpacket
		.out_endofpacket   (crosser_002_out_endofpacket),         //              .endofpacket
		.out_channel       (crosser_002_out_channel),             //              .channel
		.out_data          (crosser_002_out_data),                //              .data
		.in_empty          (1'b0),                                //   (terminated)
		.in_error          (1'b0),                                //   (terminated)
		.out_empty         (),                                    //   (terminated)
		.out_error         ()                                     //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (109),
		.BITS_PER_SYMBOL     (109),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (4),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_003 (
		.in_clk            (pcie_ip_pcie_core_clk_clk),           //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),      //  in_clk_reset.reset
		.out_clk           (clk_clk),                             //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),  // out_clk_reset.reset
		.in_ready          (width_adapter_007_src_ready),         //            in.ready
		.in_valid          (width_adapter_007_src_valid),         //              .valid
		.in_startofpacket  (width_adapter_007_src_startofpacket), //              .startofpacket
		.in_endofpacket    (width_adapter_007_src_endofpacket),   //              .endofpacket
		.in_channel        (width_adapter_007_src_channel),       //              .channel
		.in_data           (width_adapter_007_src_data),          //              .data
		.out_ready         (crosser_003_out_ready),               //           out.ready
		.out_valid         (crosser_003_out_valid),               //              .valid
		.out_startofpacket (crosser_003_out_startofpacket),       //              .startofpacket
		.out_endofpacket   (crosser_003_out_endofpacket),         //              .endofpacket
		.out_channel       (crosser_003_out_channel),             //              .channel
		.out_data          (crosser_003_out_data),                //              .data
		.in_empty          (1'b0),                                //   (terminated)
		.in_error          (1'b0),                                //   (terminated)
		.out_empty         (),                                    //   (terminated)
		.out_error         ()                                     //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (145),
		.BITS_PER_SYMBOL     (145),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (4),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_004 (
		.in_clk            (clk_clk),                             //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),  //  in_clk_reset.reset
		.out_clk           (pcie_ip_pcie_core_clk_clk),           //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),      // out_clk_reset.reset
		.in_ready          (width_adapter_010_src_ready),         //            in.ready
		.in_valid          (width_adapter_010_src_valid),         //              .valid
		.in_startofpacket  (width_adapter_010_src_startofpacket), //              .startofpacket
		.in_endofpacket    (width_adapter_010_src_endofpacket),   //              .endofpacket
		.in_channel        (width_adapter_010_src_channel),       //              .channel
		.in_data           (width_adapter_010_src_data),          //              .data
		.out_ready         (crosser_004_out_ready),               //           out.ready
		.out_valid         (crosser_004_out_valid),               //              .valid
		.out_startofpacket (crosser_004_out_startofpacket),       //              .startofpacket
		.out_endofpacket   (crosser_004_out_endofpacket),         //              .endofpacket
		.out_channel       (crosser_004_out_channel),             //              .channel
		.out_data          (crosser_004_out_data),                //              .data
		.in_empty          (1'b0),                                //   (terminated)
		.in_error          (1'b0),                                //   (terminated)
		.out_empty         (),                                    //   (terminated)
		.out_error         ()                                     //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (145),
		.BITS_PER_SYMBOL     (145),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (4),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_005 (
		.in_clk            (clk_clk),                             //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),  //  in_clk_reset.reset
		.out_clk           (pcie_ip_pcie_core_clk_clk),           //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),      // out_clk_reset.reset
		.in_ready          (width_adapter_011_src_ready),         //            in.ready
		.in_valid          (width_adapter_011_src_valid),         //              .valid
		.in_startofpacket  (width_adapter_011_src_startofpacket), //              .startofpacket
		.in_endofpacket    (width_adapter_011_src_endofpacket),   //              .endofpacket
		.in_channel        (width_adapter_011_src_channel),       //              .channel
		.in_data           (width_adapter_011_src_data),          //              .data
		.out_ready         (crosser_005_out_ready),               //           out.ready
		.out_valid         (crosser_005_out_valid),               //              .valid
		.out_startofpacket (crosser_005_out_startofpacket),       //              .startofpacket
		.out_endofpacket   (crosser_005_out_endofpacket),         //              .endofpacket
		.out_channel       (crosser_005_out_channel),             //              .channel
		.out_data          (crosser_005_out_data),                //              .data
		.in_empty          (1'b0),                                //   (terminated)
		.in_error          (1'b0),                                //   (terminated)
		.out_empty         (),                                    //   (terminated)
		.out_error         ()                                     //   (terminated)
	);

	amm_master_qsys_with_pcie_irq_mapper irq_mapper (
		.clk           (pcie_ip_pcie_core_clk_clk),      //       clk.clk
		.reset         (~pcie_ip_pcie_core_reset_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (pcie_ip_rxm_irq_irq)             //    sender.irq
	);

endmodule
