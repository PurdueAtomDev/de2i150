// amm_master_qsys_custom_with_bfm.v

// Generated using ACDS version 13.0sp1 232 at 2015.02.16.16:52:21

`timescale 1 ps / 1 ps
module amm_master_qsys_custom_with_bfm (
		input  wire        clk_clk,                            //                   clk.clk
		input  wire        reset_reset_n,                      //                 reset.reset_n
		input  wire        custom_module_conduit_rdwr_cntl,    // custom_module_conduit.rdwr_cntl
		input  wire        custom_module_conduit_n_action,     //                      .n_action
		input  wire        custom_module_conduit_add_data_sel, //                      .add_data_sel
		input  wire [25:0] custom_module_conduit_rdwr_address  //                      .rdwr_address
	);

	wire         custom_module_0_avalon_master_waitrequest;                                        // custom_module_0_avalon_master_translator:av_waitrequest -> custom_module_0:master_waitrequest
	wire  [31:0] custom_module_0_avalon_master_writedata;                                          // custom_module_0:master_writedata -> custom_module_0_avalon_master_translator:av_writedata
	wire  [25:0] custom_module_0_avalon_master_address;                                            // custom_module_0:master_address -> custom_module_0_avalon_master_translator:av_address
	wire         custom_module_0_avalon_master_write;                                              // custom_module_0:master_write -> custom_module_0_avalon_master_translator:av_write
	wire         custom_module_0_avalon_master_read;                                               // custom_module_0:master_read -> custom_module_0_avalon_master_translator:av_read
	wire  [31:0] custom_module_0_avalon_master_readdata;                                           // custom_module_0_avalon_master_translator:av_readdata -> custom_module_0:master_readdata
	wire         custom_module_0_avalon_master_readdatavalid;                                      // custom_module_0_avalon_master_translator:av_readdatavalid -> custom_module_0:master_readdatavalid
	wire         custom_module_0_avalon_master_translator_avalon_universal_master_0_waitrequest;   // mm_slave_bfm_0_s0_translator:uav_waitrequest -> custom_module_0_avalon_master_translator:uav_waitrequest
	wire   [2:0] custom_module_0_avalon_master_translator_avalon_universal_master_0_burstcount;    // custom_module_0_avalon_master_translator:uav_burstcount -> mm_slave_bfm_0_s0_translator:uav_burstcount
	wire  [31:0] custom_module_0_avalon_master_translator_avalon_universal_master_0_writedata;     // custom_module_0_avalon_master_translator:uav_writedata -> mm_slave_bfm_0_s0_translator:uav_writedata
	wire  [25:0] custom_module_0_avalon_master_translator_avalon_universal_master_0_address;       // custom_module_0_avalon_master_translator:uav_address -> mm_slave_bfm_0_s0_translator:uav_address
	wire         custom_module_0_avalon_master_translator_avalon_universal_master_0_lock;          // custom_module_0_avalon_master_translator:uav_lock -> mm_slave_bfm_0_s0_translator:uav_lock
	wire         custom_module_0_avalon_master_translator_avalon_universal_master_0_write;         // custom_module_0_avalon_master_translator:uav_write -> mm_slave_bfm_0_s0_translator:uav_write
	wire         custom_module_0_avalon_master_translator_avalon_universal_master_0_read;          // custom_module_0_avalon_master_translator:uav_read -> mm_slave_bfm_0_s0_translator:uav_read
	wire  [31:0] custom_module_0_avalon_master_translator_avalon_universal_master_0_readdata;      // mm_slave_bfm_0_s0_translator:uav_readdata -> custom_module_0_avalon_master_translator:uav_readdata
	wire         custom_module_0_avalon_master_translator_avalon_universal_master_0_debugaccess;   // custom_module_0_avalon_master_translator:uav_debugaccess -> mm_slave_bfm_0_s0_translator:uav_debugaccess
	wire   [3:0] custom_module_0_avalon_master_translator_avalon_universal_master_0_byteenable;    // custom_module_0_avalon_master_translator:uav_byteenable -> mm_slave_bfm_0_s0_translator:uav_byteenable
	wire         custom_module_0_avalon_master_translator_avalon_universal_master_0_readdatavalid; // mm_slave_bfm_0_s0_translator:uav_readdatavalid -> custom_module_0_avalon_master_translator:uav_readdatavalid
	wire         mm_slave_bfm_0_s0_translator_avalon_anti_slave_0_waitrequest;                     // mm_slave_bfm_0:avs_waitrequest -> mm_slave_bfm_0_s0_translator:av_waitrequest
	wire  [31:0] mm_slave_bfm_0_s0_translator_avalon_anti_slave_0_writedata;                       // mm_slave_bfm_0_s0_translator:av_writedata -> mm_slave_bfm_0:avs_writedata
	wire  [23:0] mm_slave_bfm_0_s0_translator_avalon_anti_slave_0_address;                         // mm_slave_bfm_0_s0_translator:av_address -> mm_slave_bfm_0:avs_address
	wire         mm_slave_bfm_0_s0_translator_avalon_anti_slave_0_write;                           // mm_slave_bfm_0_s0_translator:av_write -> mm_slave_bfm_0:avs_write
	wire         mm_slave_bfm_0_s0_translator_avalon_anti_slave_0_read;                            // mm_slave_bfm_0_s0_translator:av_read -> mm_slave_bfm_0:avs_read
	wire  [31:0] mm_slave_bfm_0_s0_translator_avalon_anti_slave_0_readdata;                        // mm_slave_bfm_0:avs_readdata -> mm_slave_bfm_0_s0_translator:av_readdata
	wire         mm_slave_bfm_0_s0_translator_avalon_anti_slave_0_readdatavalid;                   // mm_slave_bfm_0:avs_readdatavalid -> mm_slave_bfm_0_s0_translator:av_readdatavalid
	wire         mm_master_bfm_0_m0_waitrequest;                                                   // mm_master_bfm_0_m0_translator:av_waitrequest -> mm_master_bfm_0:avm_waitrequest
	wire  [31:0] mm_master_bfm_0_m0_writedata;                                                     // mm_master_bfm_0:avm_writedata -> mm_master_bfm_0_m0_translator:av_writedata
	wire  [31:0] mm_master_bfm_0_m0_address;                                                       // mm_master_bfm_0:avm_address -> mm_master_bfm_0_m0_translator:av_address
	wire         mm_master_bfm_0_m0_write;                                                         // mm_master_bfm_0:avm_write -> mm_master_bfm_0_m0_translator:av_write
	wire         mm_master_bfm_0_m0_read;                                                          // mm_master_bfm_0:avm_read -> mm_master_bfm_0_m0_translator:av_read
	wire  [31:0] mm_master_bfm_0_m0_readdata;                                                      // mm_master_bfm_0_m0_translator:av_readdata -> mm_master_bfm_0:avm_readdata
	wire         mm_master_bfm_0_m0_readdatavalid;                                                 // mm_master_bfm_0_m0_translator:av_readdatavalid -> mm_master_bfm_0:avm_readdatavalid
	wire         mm_master_bfm_0_m0_translator_avalon_universal_master_0_waitrequest;              // custom_module_0_avalon_slave_translator:uav_waitrequest -> mm_master_bfm_0_m0_translator:uav_waitrequest
	wire   [2:0] mm_master_bfm_0_m0_translator_avalon_universal_master_0_burstcount;               // mm_master_bfm_0_m0_translator:uav_burstcount -> custom_module_0_avalon_slave_translator:uav_burstcount
	wire  [31:0] mm_master_bfm_0_m0_translator_avalon_universal_master_0_writedata;                // mm_master_bfm_0_m0_translator:uav_writedata -> custom_module_0_avalon_slave_translator:uav_writedata
	wire  [31:0] mm_master_bfm_0_m0_translator_avalon_universal_master_0_address;                  // mm_master_bfm_0_m0_translator:uav_address -> custom_module_0_avalon_slave_translator:uav_address
	wire         mm_master_bfm_0_m0_translator_avalon_universal_master_0_lock;                     // mm_master_bfm_0_m0_translator:uav_lock -> custom_module_0_avalon_slave_translator:uav_lock
	wire         mm_master_bfm_0_m0_translator_avalon_universal_master_0_write;                    // mm_master_bfm_0_m0_translator:uav_write -> custom_module_0_avalon_slave_translator:uav_write
	wire         mm_master_bfm_0_m0_translator_avalon_universal_master_0_read;                     // mm_master_bfm_0_m0_translator:uav_read -> custom_module_0_avalon_slave_translator:uav_read
	wire  [31:0] mm_master_bfm_0_m0_translator_avalon_universal_master_0_readdata;                 // custom_module_0_avalon_slave_translator:uav_readdata -> mm_master_bfm_0_m0_translator:uav_readdata
	wire         mm_master_bfm_0_m0_translator_avalon_universal_master_0_debugaccess;              // mm_master_bfm_0_m0_translator:uav_debugaccess -> custom_module_0_avalon_slave_translator:uav_debugaccess
	wire   [3:0] mm_master_bfm_0_m0_translator_avalon_universal_master_0_byteenable;               // mm_master_bfm_0_m0_translator:uav_byteenable -> custom_module_0_avalon_slave_translator:uav_byteenable
	wire         mm_master_bfm_0_m0_translator_avalon_universal_master_0_readdatavalid;            // custom_module_0_avalon_slave_translator:uav_readdatavalid -> mm_master_bfm_0_m0_translator:uav_readdatavalid
	wire  [31:0] custom_module_0_avalon_slave_translator_avalon_anti_slave_0_writedata;            // custom_module_0_avalon_slave_translator:av_writedata -> custom_module_0:slave_writedata
	wire   [2:0] custom_module_0_avalon_slave_translator_avalon_anti_slave_0_address;              // custom_module_0_avalon_slave_translator:av_address -> custom_module_0:slave_address
	wire         custom_module_0_avalon_slave_translator_avalon_anti_slave_0_chipselect;           // custom_module_0_avalon_slave_translator:av_chipselect -> custom_module_0:slave_chipselect
	wire         custom_module_0_avalon_slave_translator_avalon_anti_slave_0_write;                // custom_module_0_avalon_slave_translator:av_write -> custom_module_0:slave_write
	wire         custom_module_0_avalon_slave_translator_avalon_anti_slave_0_read;                 // custom_module_0_avalon_slave_translator:av_read -> custom_module_0:slave_read
	wire  [31:0] custom_module_0_avalon_slave_translator_avalon_anti_slave_0_readdata;             // custom_module_0:slave_readdata -> custom_module_0_avalon_slave_translator:av_readdata
	wire         rst_controller_reset_out_reset;                                                   // rst_controller:reset_out -> [custom_module_0:reset, custom_module_0_avalon_master_translator:reset, custom_module_0_avalon_slave_translator:reset, mm_master_bfm_0:reset, mm_master_bfm_0_m0_translator:reset, mm_slave_bfm_0:reset, mm_slave_bfm_0_s0_translator:reset]

	altera_avalon_mm_master_bfm #(
		.AV_ADDRESS_W               (32),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (4),
		.AV_BURSTCOUNT_W            (1),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (0),
		.USE_BURSTCOUNT             (0),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (1),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_BURST_LINEWRAP          (0),
		.AV_BURST_BNDR_ONLY         (0),
		.AV_MAX_PENDING_READS       (0),
		.AV_FIX_READ_LATENCY        (1),
		.AV_READ_WAIT_TIME          (1),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (1),
		.AV_REGISTERINCOMINGSIGNALS (1),
		.VHDL_ID                    (0)
	) mm_master_bfm_0 (
		.clk                      (clk_clk),                          //       clk.clk
		.reset                    (rst_controller_reset_out_reset),   // clk_reset.reset
		.avm_address              (mm_master_bfm_0_m0_address),       //        m0.address
		.avm_readdata             (mm_master_bfm_0_m0_readdata),      //          .readdata
		.avm_writedata            (mm_master_bfm_0_m0_writedata),     //          .writedata
		.avm_waitrequest          (mm_master_bfm_0_m0_waitrequest),   //          .waitrequest
		.avm_write                (mm_master_bfm_0_m0_write),         //          .write
		.avm_read                 (mm_master_bfm_0_m0_read),          //          .read
		.avm_readdatavalid        (mm_master_bfm_0_m0_readdatavalid), //          .readdatavalid
		.avm_burstcount           (),                                 // (terminated)
		.avm_begintransfer        (),                                 // (terminated)
		.avm_beginbursttransfer   (),                                 // (terminated)
		.avm_byteenable           (),                                 // (terminated)
		.avm_arbiterlock          (),                                 // (terminated)
		.avm_lock                 (),                                 // (terminated)
		.avm_debugaccess          (),                                 // (terminated)
		.avm_transactionid        (),                                 // (terminated)
		.avm_readresponse         (8'b00000000),                      // (terminated)
		.avm_readid               (8'b00000000),                      // (terminated)
		.avm_writeresponserequest (),                                 // (terminated)
		.avm_writeresponse        (8'b00000000),                      // (terminated)
		.avm_writeresponsevalid   (1'b0),                             // (terminated)
		.avm_writeid              (8'b00000000),                      // (terminated)
		.avm_clken                ()                                  // (terminated)
	);

	altera_avalon_mm_slave_bfm #(
		.AV_ADDRESS_W               (24),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (4),
		.AV_BURSTCOUNT_W            (3),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (0),
		.USE_BURSTCOUNT             (0),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (1),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_BURST_LINEWRAP          (0),
		.AV_BURST_BNDR_ONLY         (0),
		.AV_MAX_PENDING_READS       (1),
		.AV_FIX_READ_LATENCY        (0),
		.AV_READ_WAIT_TIME          (1),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (0)
	) mm_slave_bfm_0 (
		.clk                      (clk_clk),                                                        //       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                 // clk_reset.reset
		.avs_writedata            (mm_slave_bfm_0_s0_translator_avalon_anti_slave_0_writedata),     //        s0.writedata
		.avs_readdata             (mm_slave_bfm_0_s0_translator_avalon_anti_slave_0_readdata),      //          .readdata
		.avs_address              (mm_slave_bfm_0_s0_translator_avalon_anti_slave_0_address),       //          .address
		.avs_waitrequest          (mm_slave_bfm_0_s0_translator_avalon_anti_slave_0_waitrequest),   //          .waitrequest
		.avs_write                (mm_slave_bfm_0_s0_translator_avalon_anti_slave_0_write),         //          .write
		.avs_read                 (mm_slave_bfm_0_s0_translator_avalon_anti_slave_0_read),          //          .read
		.avs_readdatavalid        (mm_slave_bfm_0_s0_translator_avalon_anti_slave_0_readdatavalid), //          .readdatavalid
		.avs_begintransfer        (1'b0),                                                           // (terminated)
		.avs_beginbursttransfer   (1'b0),                                                           // (terminated)
		.avs_burstcount           (3'b001),                                                         // (terminated)
		.avs_byteenable           (4'b1111),                                                        // (terminated)
		.avs_arbiterlock          (1'b0),                                                           // (terminated)
		.avs_lock                 (1'b0),                                                           // (terminated)
		.avs_debugaccess          (1'b0),                                                           // (terminated)
		.avs_transactionid        (8'b00000000),                                                    // (terminated)
		.avs_readresponse         (),                                                               // (terminated)
		.avs_readid               (),                                                               // (terminated)
		.avs_writeresponserequest (1'b0),                                                           // (terminated)
		.avs_writeresponse        (),                                                               // (terminated)
		.avs_writeresponsevalid   (),                                                               // (terminated)
		.avs_writeid              (),                                                               // (terminated)
		.avs_clken                (1'b1)                                                            // (terminated)
	);

	custom_slave #(
		.MASTER_ADDRESSWIDTH (26),
		.SLAVE_ADDRESSWIDTH  (3),
		.DATAWIDTH           (32),
		.NUMREGS             (8),
		.REGWIDTH            (32)
	) custom_module_0 (
		.clk                  (clk_clk),                                                                //         clock.clk
		.reset_n                (~rst_controller_reset_out_reset),                                        //         reset.reset_n
		.master_address       (custom_module_0_avalon_master_address),                                  // avalon_master.address
		.master_writedata     (custom_module_0_avalon_master_writedata),                                //              .writedata
		.master_write         (custom_module_0_avalon_master_write),                                    //              .write
		.master_read          (custom_module_0_avalon_master_read),                                     //              .read
		.master_readdata      (custom_module_0_avalon_master_readdata),                                 //              .readdata
		.master_readdatavalid (custom_module_0_avalon_master_readdatavalid),                            //              .readdatavalid
		.master_waitrequest   (custom_module_0_avalon_master_waitrequest),                              //              .waitrequest
		.slave_readdata       (custom_module_0_avalon_slave_translator_avalon_anti_slave_0_readdata),   //  avalon_slave.readdata
		.slave_chipselect     (custom_module_0_avalon_slave_translator_avalon_anti_slave_0_chipselect), //              .chipselect
		.slave_read           (custom_module_0_avalon_slave_translator_avalon_anti_slave_0_read),       //              .read
		.slave_write          (custom_module_0_avalon_slave_translator_avalon_anti_slave_0_write),      //              .write
		.slave_writedata      (custom_module_0_avalon_slave_translator_avalon_anti_slave_0_writedata),  //              .writedata
		.slave_address        (custom_module_0_avalon_slave_translator_avalon_anti_slave_0_address),    //              .address
		.rdwr_cntl            (custom_module_conduit_rdwr_cntl),                                        //   conduit_end.export
		.n_action             (custom_module_conduit_n_action),                                         //              .export
		.add_data_sel         (custom_module_conduit_add_data_sel),                                     //              .export
		.rdwr_address         (custom_module_conduit_rdwr_address)                                      //              .export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (26),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (26),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) custom_module_0_avalon_master_translator (
		.clk                      (clk_clk),                                                                          //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                   //                     reset.reset
		.uav_address              (custom_module_0_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (custom_module_0_avalon_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (custom_module_0_avalon_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (custom_module_0_avalon_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (custom_module_0_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (custom_module_0_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (custom_module_0_avalon_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (custom_module_0_avalon_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (custom_module_0_avalon_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (custom_module_0_avalon_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (custom_module_0_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (custom_module_0_avalon_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (custom_module_0_avalon_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (custom_module_0_avalon_master_read),                                               //                          .read
		.av_readdata              (custom_module_0_avalon_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (custom_module_0_avalon_master_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (custom_module_0_avalon_master_write),                                              //                          .write
		.av_writedata             (custom_module_0_avalon_master_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                             //               (terminated)
		.av_byteenable            (4'b1111),                                                                          //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                             //               (terminated)
		.av_begintransfer         (1'b0),                                                                             //               (terminated)
		.av_chipselect            (1'b0),                                                                             //               (terminated)
		.av_lock                  (1'b0),                                                                             //               (terminated)
		.av_debugaccess           (1'b0),                                                                             //               (terminated)
		.uav_clken                (),                                                                                 //               (terminated)
		.av_clken                 (1'b1),                                                                             //               (terminated)
		.uav_response             (2'b00),                                                                            //               (terminated)
		.av_response              (),                                                                                 //               (terminated)
		.uav_writeresponserequest (),                                                                                 //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                             //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                             //               (terminated)
		.av_writeresponsevalid    ()                                                                                  //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (24),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) mm_slave_bfm_0_s0_translator (
		.clk                      (clk_clk),                                                                          //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                   //                    reset.reset
		.uav_address              (custom_module_0_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (custom_module_0_avalon_master_translator_avalon_universal_master_0_burstcount),    //                         .burstcount
		.uav_read                 (custom_module_0_avalon_master_translator_avalon_universal_master_0_read),          //                         .read
		.uav_write                (custom_module_0_avalon_master_translator_avalon_universal_master_0_write),         //                         .write
		.uav_waitrequest          (custom_module_0_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (custom_module_0_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (custom_module_0_avalon_master_translator_avalon_universal_master_0_byteenable),    //                         .byteenable
		.uav_readdata             (custom_module_0_avalon_master_translator_avalon_universal_master_0_readdata),      //                         .readdata
		.uav_writedata            (custom_module_0_avalon_master_translator_avalon_universal_master_0_writedata),     //                         .writedata
		.uav_lock                 (custom_module_0_avalon_master_translator_avalon_universal_master_0_lock),          //                         .lock
		.uav_debugaccess          (custom_module_0_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                         .debugaccess
		.av_address               (mm_slave_bfm_0_s0_translator_avalon_anti_slave_0_address),                         //      avalon_anti_slave_0.address
		.av_write                 (mm_slave_bfm_0_s0_translator_avalon_anti_slave_0_write),                           //                         .write
		.av_read                  (mm_slave_bfm_0_s0_translator_avalon_anti_slave_0_read),                            //                         .read
		.av_readdata              (mm_slave_bfm_0_s0_translator_avalon_anti_slave_0_readdata),                        //                         .readdata
		.av_writedata             (mm_slave_bfm_0_s0_translator_avalon_anti_slave_0_writedata),                       //                         .writedata
		.av_readdatavalid         (mm_slave_bfm_0_s0_translator_avalon_anti_slave_0_readdatavalid),                   //                         .readdatavalid
		.av_waitrequest           (mm_slave_bfm_0_s0_translator_avalon_anti_slave_0_waitrequest),                     //                         .waitrequest
		.av_begintransfer         (),                                                                                 //              (terminated)
		.av_beginbursttransfer    (),                                                                                 //              (terminated)
		.av_burstcount            (),                                                                                 //              (terminated)
		.av_byteenable            (),                                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                                 //              (terminated)
		.av_lock                  (),                                                                                 //              (terminated)
		.av_chipselect            (),                                                                                 //              (terminated)
		.av_clken                 (),                                                                                 //              (terminated)
		.uav_clken                (1'b0),                                                                             //              (terminated)
		.av_debugaccess           (),                                                                                 //              (terminated)
		.av_outputenable          (),                                                                                 //              (terminated)
		.uav_response             (),                                                                                 //              (terminated)
		.av_response              (2'b00),                                                                            //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                             //              (terminated)
		.uav_writeresponsevalid   (),                                                                                 //              (terminated)
		.av_writeresponserequest  (),                                                                                 //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                              //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) mm_master_bfm_0_m0_translator (
		.clk                      (clk_clk),                                                               //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                     reset.reset
		.uav_address              (mm_master_bfm_0_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (mm_master_bfm_0_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (mm_master_bfm_0_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (mm_master_bfm_0_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (mm_master_bfm_0_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (mm_master_bfm_0_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (mm_master_bfm_0_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (mm_master_bfm_0_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (mm_master_bfm_0_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (mm_master_bfm_0_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (mm_master_bfm_0_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (mm_master_bfm_0_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (mm_master_bfm_0_m0_waitrequest),                                        //                          .waitrequest
		.av_read                  (mm_master_bfm_0_m0_read),                                               //                          .read
		.av_readdata              (mm_master_bfm_0_m0_readdata),                                           //                          .readdata
		.av_readdatavalid         (mm_master_bfm_0_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (mm_master_bfm_0_m0_write),                                              //                          .write
		.av_writedata             (mm_master_bfm_0_m0_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                  //               (terminated)
		.av_byteenable            (4'b1111),                                                               //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                  //               (terminated)
		.av_begintransfer         (1'b0),                                                                  //               (terminated)
		.av_chipselect            (1'b0),                                                                  //               (terminated)
		.av_lock                  (1'b0),                                                                  //               (terminated)
		.av_debugaccess           (1'b0),                                                                  //               (terminated)
		.uav_clken                (),                                                                      //               (terminated)
		.av_clken                 (1'b1),                                                                  //               (terminated)
		.uav_response             (2'b00),                                                                 //               (terminated)
		.av_response              (),                                                                      //               (terminated)
		.uav_writeresponserequest (),                                                                      //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                  //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                  //               (terminated)
		.av_writeresponsevalid    ()                                                                       //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) custom_module_0_avalon_slave_translator (
		.clk                      (clk_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                         //                    reset.reset
		.uav_address              (mm_master_bfm_0_m0_translator_avalon_universal_master_0_address),        // avalon_universal_slave_0.address
		.uav_burstcount           (mm_master_bfm_0_m0_translator_avalon_universal_master_0_burstcount),     //                         .burstcount
		.uav_read                 (mm_master_bfm_0_m0_translator_avalon_universal_master_0_read),           //                         .read
		.uav_write                (mm_master_bfm_0_m0_translator_avalon_universal_master_0_write),          //                         .write
		.uav_waitrequest          (mm_master_bfm_0_m0_translator_avalon_universal_master_0_waitrequest),    //                         .waitrequest
		.uav_readdatavalid        (mm_master_bfm_0_m0_translator_avalon_universal_master_0_readdatavalid),  //                         .readdatavalid
		.uav_byteenable           (mm_master_bfm_0_m0_translator_avalon_universal_master_0_byteenable),     //                         .byteenable
		.uav_readdata             (mm_master_bfm_0_m0_translator_avalon_universal_master_0_readdata),       //                         .readdata
		.uav_writedata            (mm_master_bfm_0_m0_translator_avalon_universal_master_0_writedata),      //                         .writedata
		.uav_lock                 (mm_master_bfm_0_m0_translator_avalon_universal_master_0_lock),           //                         .lock
		.uav_debugaccess          (mm_master_bfm_0_m0_translator_avalon_universal_master_0_debugaccess),    //                         .debugaccess
		.av_address               (custom_module_0_avalon_slave_translator_avalon_anti_slave_0_address),    //      avalon_anti_slave_0.address
		.av_write                 (custom_module_0_avalon_slave_translator_avalon_anti_slave_0_write),      //                         .write
		.av_read                  (custom_module_0_avalon_slave_translator_avalon_anti_slave_0_read),       //                         .read
		.av_readdata              (custom_module_0_avalon_slave_translator_avalon_anti_slave_0_readdata),   //                         .readdata
		.av_writedata             (custom_module_0_avalon_slave_translator_avalon_anti_slave_0_writedata),  //                         .writedata
		.av_chipselect            (custom_module_0_avalon_slave_translator_avalon_anti_slave_0_chipselect), //                         .chipselect
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

endmodule
